module ff_tcam_tb();
parameter BITADDR = 4;
parameter WIDTH = 10;

reg clk, rst;




endmodule
