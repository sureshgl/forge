module topModule;

slave1 u_slave1 ();

slave2 u_slave2 ();

slave3 u_slave3 ();


endmodule