`define ARB_FIFO_PKT_THRESHOLD_0_OFFSET	32'h0
`define ARB_FIFO_PKT_THRESHOLD_0_SIZE	16
`define ARB_FIFO_PKT_THRESHOLD_0_SIZE_IN_WORDS	1

`define ARB_FIFO_PKT_THRESHOLD_0_THRESH_SIZE	16
`define ARB_FIFO_PKT_THRESHOLD_0_THRESH_START_OFFSET	0
`define ARB_FIFO_PKT_THRESHOLD_0_THRESH_RANGE	[15:0]
`define ARB_FIFO_PKT_THRESHOLD_0_THRESH_RST_VALUE	16'hF0




`define PROC_PKT_THRESHOLD_0_OFFSET	32'h4
`define PROC_PKT_THRESHOLD_0_SIZE	33
`define PROC_PKT_THRESHOLD_0_SIZE_IN_WORDS	2

`define PROC_PKT_THRESHOLD_0_THRESH_SIZE	30
`define PROC_PKT_THRESHOLD_0_THRESH_START_OFFSET	0
`define PROC_PKT_THRESHOLD_0_THRESH_RANGE	[29:0]
`define PROC_PKT_THRESHOLD_0_THRESH_RST_VALUE	30'h0

`define PROC_PKT_THRESHOLD_0_THR_SIZE	3
`define PROC_PKT_THRESHOLD_0_THR_START_OFFSET	30
`define PROC_PKT_THRESHOLD_0_THR_RANGE	[32:30]
`define PROC_PKT_THRESHOLD_0_THR_RST_VALUE	16'h0FF



`define PROC_PKT_THRESHOLD_1_OFFSET	32'h6
`define PROC_PKT_THRESHOLD_1_SIZE	33
`define PROC_PKT_THRESHOLD_1_SIZE_IN_WORDS	2

`define PROC_PKT_THRESHOLD_1_THRESH_SIZE	30
`define PROC_PKT_THRESHOLD_1_THRESH_START_OFFSET	0
`define PROC_PKT_THRESHOLD_1_THRESH_RANGE	[29:0]
`define PROC_PKT_THRESHOLD_1_THRESH_RST_VALUE	30'h0

`define PROC_PKT_THRESHOLD_1_THR_SIZE	3
`define PROC_PKT_THRESHOLD_1_THR_START_OFFSET	30
`define PROC_PKT_THRESHOLD_1_THR_RANGE	[32:30]
`define PROC_PKT_THRESHOLD_1_THR_RST_VALUE	16'h0FF



`define PROC_PKT_THRESHOLD_2_OFFSET	32'h8
`define PROC_PKT_THRESHOLD_2_SIZE	33
`define PROC_PKT_THRESHOLD_2_SIZE_IN_WORDS	2

`define PROC_PKT_THRESHOLD_2_THRESH_SIZE	30
`define PROC_PKT_THRESHOLD_2_THRESH_START_OFFSET	0
`define PROC_PKT_THRESHOLD_2_THRESH_RANGE	[29:0]
`define PROC_PKT_THRESHOLD_2_THRESH_RST_VALUE	30'h0

`define PROC_PKT_THRESHOLD_2_THR_SIZE	3
`define PROC_PKT_THRESHOLD_2_THR_START_OFFSET	30
`define PROC_PKT_THRESHOLD_2_THR_RANGE	[32:30]
`define PROC_PKT_THRESHOLD_2_THR_RST_VALUE	16'h0FF




`define DUMMYREG_0_OFFSET	32'h8
`define DUMMYREG_0_SIZE	39
`define DUMMYREG_0_SIZE_IN_WORDS	2

`define DUMMYREG_0_THRESH_SIZE	39
`define DUMMYREG_0_THRESH_START_OFFSET	0
`define DUMMYREG_0_THRESH_RANGE	[38:0]
`define DUMMYREG_0_THRESH_RST_VALUE	16'hF0




`define DUMMY_REG1_0_OFFSET	32'h20
`define DUMMY_REG1_0_SIZE	65
`define DUMMY_REG1_0_SIZE_IN_WORDS	3

`define DUMMY_REG1_0_THRESH_SIZE	65
`define DUMMY_REG1_0_THRESH_START_OFFSET	0
`define DUMMY_REG1_0_THRESH_RANGE	[64:0]
`define DUMMY_REG1_0_THRESH_RST_VALUE	16'h0FF



`define DUMMY_REG1_1_OFFSET	32'h23
`define DUMMY_REG1_1_SIZE	65
`define DUMMY_REG1_1_SIZE_IN_WORDS	3

`define DUMMY_REG1_1_THRESH_SIZE	65
`define DUMMY_REG1_1_THRESH_START_OFFSET	0
`define DUMMY_REG1_1_THRESH_RANGE	[64:0]
`define DUMMY_REG1_1_THRESH_RST_VALUE	16'h0FF



`define DUMMY_REG1_2_OFFSET	32'h26
`define DUMMY_REG1_2_SIZE	65
`define DUMMY_REG1_2_SIZE_IN_WORDS	3

`define DUMMY_REG1_2_THRESH_SIZE	65
`define DUMMY_REG1_2_THRESH_START_OFFSET	0
`define DUMMY_REG1_2_THRESH_RANGE	[64:0]
`define DUMMY_REG1_2_THRESH_RST_VALUE	16'h0FF



`define DUMMY_REG1_3_OFFSET	32'h29
`define DUMMY_REG1_3_SIZE	65
`define DUMMY_REG1_3_SIZE_IN_WORDS	3

`define DUMMY_REG1_3_THRESH_SIZE	65
`define DUMMY_REG1_3_THRESH_START_OFFSET	0
`define DUMMY_REG1_3_THRESH_RANGE	[64:0]
`define DUMMY_REG1_3_THRESH_RST_VALUE	16'h0FF



`define DUMMY_REG1_4_OFFSET	32'h2c
`define DUMMY_REG1_4_SIZE	65
`define DUMMY_REG1_4_SIZE_IN_WORDS	3

`define DUMMY_REG1_4_THRESH_SIZE	65
`define DUMMY_REG1_4_THRESH_START_OFFSET	0
`define DUMMY_REG1_4_THRESH_RANGE	[64:0]
`define DUMMY_REG1_4_THRESH_RST_VALUE	16'h0FF



`define DUMMY_REG1_5_OFFSET	32'h2f
`define DUMMY_REG1_5_SIZE	65
`define DUMMY_REG1_5_SIZE_IN_WORDS	3

`define DUMMY_REG1_5_THRESH_SIZE	65
`define DUMMY_REG1_5_THRESH_START_OFFSET	0
`define DUMMY_REG1_5_THRESH_RANGE	[64:0]
`define DUMMY_REG1_5_THRESH_RST_VALUE	16'h0FF





