`ifdef __DCMDESC_VH__
`else
`define __DCMDESC_VH__

// Defines for DcmDesc

// macros for register Dcm_DeskewTableDesc
//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tsq0DeskewCount
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_RANGE                       7:0
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_MSB                           7
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_LSB                           0
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_REL_RANGE                   7:0
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_REL_MSB                       7
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_REL_LSB                       0
`define DCM_DESKEWTABLEDESC_TSQ0DESKEWCOUNT_RESET_VALUE               8'hb6

// macros with short names for field Dcm_DeskewTableDesc.tsq0DeskewCount
`define DCM_DSKWTBLDSC_TSQ0DSKWCNT_RANGE                                7:0
`define DCM_DSKWTBLDSC_TSQ0DSKWCNT_MSB                                    7
`define DCM_DSKWTBLDSC_TSQ0DSKWCNT_LSB                                    0
`define DCM_DSKWTBLDSC_TSQ0DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TSQ0DSKWCNT_RESET_VALUE                        8'hb6

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tsq1DeskewCount
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_RANGE                      15:8
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_MSB                          15
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_LSB                           8
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_REL_RANGE                  15:8
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_REL_MSB                      15
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_REL_LSB                       8
`define DCM_DESKEWTABLEDESC_TSQ1DESKEWCOUNT_RESET_VALUE               8'hb5

// macros with short names for field Dcm_DeskewTableDesc.tsq1DeskewCount
`define DCM_DSKWTBLDSC_TSQ1DSKWCNT_RANGE                               15:8
`define DCM_DSKWTBLDSC_TSQ1DSKWCNT_MSB                                   15
`define DCM_DSKWTBLDSC_TSQ1DSKWCNT_LSB                                    8
`define DCM_DSKWTBLDSC_TSQ1DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TSQ1DSKWCNT_RESET_VALUE                        8'hb5

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tsq2DeskewCount
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_RANGE                     23:16
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_MSB                          23
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_LSB                          16
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_REL_RANGE                 23:16
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_REL_MSB                      23
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_REL_LSB                      16
`define DCM_DESKEWTABLEDESC_TSQ2DESKEWCOUNT_RESET_VALUE               8'hb4

// macros with short names for field Dcm_DeskewTableDesc.tsq2DeskewCount
`define DCM_DSKWTBLDSC_TSQ2DSKWCNT_RANGE                              23:16
`define DCM_DSKWTBLDSC_TSQ2DSKWCNT_MSB                                   23
`define DCM_DSKWTBLDSC_TSQ2DSKWCNT_LSB                                   16
`define DCM_DSKWTBLDSC_TSQ2DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TSQ2DSKWCNT_RESET_VALUE                        8'hb4

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tsq3DeskewCount
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_RANGE                     31:24
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_MSB                          31
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_LSB                          24
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_REL_RANGE                 31:24
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_REL_MSB                      31
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_REL_LSB                      24
`define DCM_DESKEWTABLEDESC_TSQ3DESKEWCOUNT_RESET_VALUE               8'hb4

// macros with short names for field Dcm_DeskewTableDesc.tsq3DeskewCount
`define DCM_DSKWTBLDSC_TSQ3DSKWCNT_RANGE                              31:24
`define DCM_DSKWTBLDSC_TSQ3DSKWCNT_MSB                                   31
`define DCM_DSKWTBLDSC_TSQ3DSKWCNT_LSB                                   24
`define DCM_DSKWTBLDSC_TSQ3DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TSQ3DSKWCNT_RESET_VALUE                        8'hb4

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.plcDeskewCount
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_RANGE                      39:32
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_MSB                           39
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_LSB                           32
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_REL_RANGE                  39:32
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_REL_MSB                       39
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_REL_LSB                       32
`define DCM_DESKEWTABLEDESC_PLCDESKEWCOUNT_RESET_VALUE                8'hb3

// macros with short names for field Dcm_DeskewTableDesc.plcDeskewCount
`define DCM_DSKWTBLDSC_PLCDSKWCNT_RANGE                               39:32
`define DCM_DSKWTBLDSC_PLCDSKWCNT_MSB                                    39
`define DCM_DSKWTBLDSC_PLCDSKWCNT_LSB                                    32
`define DCM_DSKWTBLDSC_PLCDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_PLCDSKWCNT_RESET_VALUE                         8'hb3

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.nflDeskewCount
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_RANGE                      47:40
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_MSB                           47
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_LSB                           40
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_REL_RANGE                  47:40
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_REL_MSB                       47
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_REL_LSB                       40
`define DCM_DESKEWTABLEDESC_NFLDESKEWCOUNT_RESET_VALUE                8'hb2

// macros with short names for field Dcm_DeskewTableDesc.nflDeskewCount
`define DCM_DSKWTBLDSC_NFLDSKWCNT_RANGE                               47:40
`define DCM_DSKWTBLDSC_NFLDSKWCNT_MSB                                    47
`define DCM_DSKWTBLDSC_NFLDSKWCNT_LSB                                    40
`define DCM_DSKWTBLDSC_NFLDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_NFLDSKWCNT_RESET_VALUE                         8'hb2

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm11DeskewCount
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_RANGE                    55:48
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_MSB                         55
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_LSB                         48
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_REL_RANGE                55:48
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_REL_MSB                     55
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_REL_LSB                     48
`define DCM_DESKEWTABLEDESC_DMM11DESKEWCOUNT_RESET_VALUE              8'hae

// macros with short names for field Dcm_DeskewTableDesc.dmm11DeskewCount
`define DCM_DSKWTBLDSC_DMM11DSKWCNT_RANGE                             55:48
`define DCM_DSKWTBLDSC_DMM11DSKWCNT_MSB                                  55
`define DCM_DSKWTBLDSC_DMM11DSKWCNT_LSB                                  48
`define DCM_DSKWTBLDSC_DMM11DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM11DSKWCNT_RESET_VALUE                       8'hae

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase0DeskewCount
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_RANGE                     63:56
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_MSB                          63
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_LSB                          56
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_REL_RANGE                 63:56
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_REL_MSB                      63
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_REL_LSB                      56
`define DCM_DESKEWTABLEDESC_ASE0DESKEWCOUNT_RESET_VALUE               8'had

// macros with short names for field Dcm_DeskewTableDesc.ase0DeskewCount
`define DCM_DSKWTBLDSC_AS0DSKWCNT_RANGE                               63:56
`define DCM_DSKWTBLDSC_AS0DSKWCNT_MSB                                    63
`define DCM_DSKWTBLDSC_AS0DSKWCNT_LSB                                    56
`define DCM_DSKWTBLDSC_AS0DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS0DSKWCNT_RESET_VALUE                         8'had

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase1DeskewCount
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_RANGE                     71:64
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_MSB                          71
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_LSB                          64
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_REL_RANGE                 71:64
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_REL_MSB                      71
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_REL_LSB                      64
`define DCM_DESKEWTABLEDESC_ASE1DESKEWCOUNT_RESET_VALUE               8'hab

// macros with short names for field Dcm_DeskewTableDesc.ase1DeskewCount
`define DCM_DSKWTBLDSC_AS1DSKWCNT_RANGE                               71:64
`define DCM_DSKWTBLDSC_AS1DSKWCNT_MSB                                    71
`define DCM_DSKWTBLDSC_AS1DSKWCNT_LSB                                    64
`define DCM_DSKWTBLDSC_AS1DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS1DSKWCNT_RESET_VALUE                         8'hab

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase2DeskewCount
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_RANGE                     79:72
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_MSB                          79
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_LSB                          72
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_REL_RANGE                 79:72
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_REL_MSB                      79
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_REL_LSB                      72
`define DCM_DESKEWTABLEDESC_ASE2DESKEWCOUNT_RESET_VALUE               8'ha9

// macros with short names for field Dcm_DeskewTableDesc.ase2DeskewCount
`define DCM_DSKWTBLDSC_AS2DSKWCNT_RANGE                               79:72
`define DCM_DSKWTBLDSC_AS2DSKWCNT_MSB                                    79
`define DCM_DSKWTBLDSC_AS2DSKWCNT_LSB                                    72
`define DCM_DSKWTBLDSC_AS2DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS2DSKWCNT_RESET_VALUE                         8'ha9

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase3DeskewCount
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_RANGE                     87:80
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_MSB                          87
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_LSB                          80
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_REL_RANGE                 87:80
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_REL_MSB                      87
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_REL_LSB                      80
`define DCM_DESKEWTABLEDESC_ASE3DESKEWCOUNT_RESET_VALUE               8'ha7

// macros with short names for field Dcm_DeskewTableDesc.ase3DeskewCount
`define DCM_DSKWTBLDSC_AS3DSKWCNT_RANGE                               87:80
`define DCM_DSKWTBLDSC_AS3DSKWCNT_MSB                                    87
`define DCM_DSKWTBLDSC_AS3DSKWCNT_LSB                                    80
`define DCM_DSKWTBLDSC_AS3DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS3DSKWCNT_RESET_VALUE                         8'ha7

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase4DeskewCount
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_RANGE                     95:88
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_MSB                          95
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_LSB                          88
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_REL_RANGE                 95:88
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_REL_MSB                      95
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_REL_LSB                      88
`define DCM_DESKEWTABLEDESC_ASE4DESKEWCOUNT_RESET_VALUE               8'ha5

// macros with short names for field Dcm_DeskewTableDesc.ase4DeskewCount
`define DCM_DSKWTBLDSC_AS4DSKWCNT_RANGE                               95:88
`define DCM_DSKWTBLDSC_AS4DSKWCNT_MSB                                    95
`define DCM_DSKWTBLDSC_AS4DSKWCNT_LSB                                    88
`define DCM_DSKWTBLDSC_AS4DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS4DSKWCNT_RESET_VALUE                         8'ha5

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase5DeskewCount
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_RANGE                    103:96
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_MSB                         103
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_LSB                          96
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_REL_RANGE                103:96
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_REL_MSB                     103
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_REL_LSB                      96
`define DCM_DESKEWTABLEDESC_ASE5DESKEWCOUNT_RESET_VALUE               8'ha3

// macros with short names for field Dcm_DeskewTableDesc.ase5DeskewCount
`define DCM_DSKWTBLDSC_AS5DSKWCNT_RANGE                              103:96
`define DCM_DSKWTBLDSC_AS5DSKWCNT_MSB                                   103
`define DCM_DSKWTBLDSC_AS5DSKWCNT_LSB                                    96
`define DCM_DSKWTBLDSC_AS5DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS5DSKWCNT_RESET_VALUE                         8'ha3

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase6DeskewCount
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_RANGE                   111:104
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_MSB                         111
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_LSB                         104
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_REL_RANGE               111:104
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_REL_MSB                     111
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_REL_LSB                     104
`define DCM_DESKEWTABLEDESC_ASE6DESKEWCOUNT_RESET_VALUE               8'ha3

// macros with short names for field Dcm_DeskewTableDesc.ase6DeskewCount
`define DCM_DSKWTBLDSC_AS6DSKWCNT_RANGE                             111:104
`define DCM_DSKWTBLDSC_AS6DSKWCNT_MSB                                   111
`define DCM_DSKWTBLDSC_AS6DSKWCNT_LSB                                   104
`define DCM_DSKWTBLDSC_AS6DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS6DSKWCNT_RESET_VALUE                         8'ha3

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ase7DeskewCount
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_RANGE                   119:112
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_MSB                         119
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_LSB                         112
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_REL_RANGE               119:112
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_REL_MSB                     119
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_REL_LSB                     112
`define DCM_DESKEWTABLEDESC_ASE7DESKEWCOUNT_RESET_VALUE               8'ha3

// macros with short names for field Dcm_DeskewTableDesc.ase7DeskewCount
`define DCM_DSKWTBLDSC_AS7DSKWCNT_RANGE                             119:112
`define DCM_DSKWTBLDSC_AS7DSKWCNT_MSB                                   119
`define DCM_DSKWTBLDSC_AS7DSKWCNT_LSB                                   112
`define DCM_DSKWTBLDSC_AS7DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AS7DSKWCNT_RESET_VALUE                         8'ha3

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.taq0DeskewCount
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_RANGE                   127:120
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_MSB                         127
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_LSB                         120
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_REL_RANGE               127:120
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_REL_MSB                     127
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_REL_LSB                     120
`define DCM_DESKEWTABLEDESC_TAQ0DESKEWCOUNT_RESET_VALUE               8'ha1

// macros with short names for field Dcm_DeskewTableDesc.taq0DeskewCount
`define DCM_DSKWTBLDSC_TQ0DSKWCNT_RANGE                             127:120
`define DCM_DSKWTBLDSC_TQ0DSKWCNT_MSB                                   127
`define DCM_DSKWTBLDSC_TQ0DSKWCNT_LSB                                   120
`define DCM_DSKWTBLDSC_TQ0DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_TQ0DSKWCNT_RESET_VALUE                         8'ha1

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.taq1DeskewCount
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_RANGE                   135:128
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_MSB                         135
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_LSB                         128
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_REL_RANGE               135:128
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_REL_MSB                     135
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_REL_LSB                     128
`define DCM_DESKEWTABLEDESC_TAQ1DESKEWCOUNT_RESET_VALUE               8'h9f

// macros with short names for field Dcm_DeskewTableDesc.taq1DeskewCount
`define DCM_DSKWTBLDSC_TQ1DSKWCNT_RANGE                             135:128
`define DCM_DSKWTBLDSC_TQ1DSKWCNT_MSB                                   135
`define DCM_DSKWTBLDSC_TQ1DSKWCNT_LSB                                   128
`define DCM_DSKWTBLDSC_TQ1DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_TQ1DSKWCNT_RESET_VALUE                         8'h9f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.taq2DeskewCount
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_RANGE                   143:136
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_MSB                         143
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_LSB                         136
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_REL_RANGE               143:136
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_REL_MSB                     143
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_REL_LSB                     136
`define DCM_DESKEWTABLEDESC_TAQ2DESKEWCOUNT_RESET_VALUE               8'h9d

// macros with short names for field Dcm_DeskewTableDesc.taq2DeskewCount
`define DCM_DSKWTBLDSC_TQ2DSKWCNT_RANGE                             143:136
`define DCM_DSKWTBLDSC_TQ2DSKWCNT_MSB                                   143
`define DCM_DSKWTBLDSC_TQ2DSKWCNT_LSB                                   136
`define DCM_DSKWTBLDSC_TQ2DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_TQ2DSKWCNT_RESET_VALUE                         8'h9d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.taq3DeskewCount
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_RANGE                   151:144
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_MSB                         151
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_LSB                         144
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_REL_RANGE               151:144
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_REL_MSB                     151
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_REL_LSB                     144
`define DCM_DESKEWTABLEDESC_TAQ3DESKEWCOUNT_RESET_VALUE               8'h9b

// macros with short names for field Dcm_DeskewTableDesc.taq3DeskewCount
`define DCM_DSKWTBLDSC_TQ3DSKWCNT_RANGE                             151:144
`define DCM_DSKWTBLDSC_TQ3DSKWCNT_MSB                                   151
`define DCM_DSKWTBLDSC_TQ3DSKWCNT_LSB                                   144
`define DCM_DSKWTBLDSC_TQ3DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_TQ3DSKWCNT_RESET_VALUE                         8'h9b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.taq4DeskewCount
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_RANGE                   159:152
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_MSB                         159
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_LSB                         152
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_REL_RANGE               159:152
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_REL_MSB                     159
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_REL_LSB                     152
`define DCM_DESKEWTABLEDESC_TAQ4DESKEWCOUNT_RESET_VALUE               8'h99

// macros with short names for field Dcm_DeskewTableDesc.taq4DeskewCount
`define DCM_DSKWTBLDSC_TQ4DSKWCNT_RANGE                             159:152
`define DCM_DSKWTBLDSC_TQ4DSKWCNT_MSB                                   159
`define DCM_DSKWTBLDSC_TQ4DSKWCNT_LSB                                   152
`define DCM_DSKWTBLDSC_TQ4DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_TQ4DSKWCNT_RESET_VALUE                         8'h99

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.taq5DeskewCount
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_RANGE                   167:160
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_MSB                         167
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_LSB                         160
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_REL_RANGE               167:160
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_REL_MSB                     167
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_REL_LSB                     160
`define DCM_DESKEWTABLEDESC_TAQ5DESKEWCOUNT_RESET_VALUE               8'h97

// macros with short names for field Dcm_DeskewTableDesc.taq5DeskewCount
`define DCM_DSKWTBLDSC_TQ5DSKWCNT_RANGE                             167:160
`define DCM_DSKWTBLDSC_TQ5DSKWCNT_MSB                                   167
`define DCM_DSKWTBLDSC_TQ5DSKWCNT_LSB                                   160
`define DCM_DSKWTBLDSC_TQ5DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_TQ5DSKWCNT_RESET_VALUE                         8'h97

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.taq6DeskewCount
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_RANGE                   175:168
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_MSB                         175
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_LSB                         168
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_REL_RANGE               175:168
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_REL_MSB                     175
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_REL_LSB                     168
`define DCM_DESKEWTABLEDESC_TAQ6DESKEWCOUNT_RESET_VALUE               8'h95

// macros with short names for field Dcm_DeskewTableDesc.taq6DeskewCount
`define DCM_DSKWTBLDSC_TQ6DSKWCNT_RANGE                             175:168
`define DCM_DSKWTBLDSC_TQ6DSKWCNT_MSB                                   175
`define DCM_DSKWTBLDSC_TQ6DSKWCNT_LSB                                   168
`define DCM_DSKWTBLDSC_TQ6DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_TQ6DSKWCNT_RESET_VALUE                         8'h95

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tlq0DeskewCount
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_RANGE                   183:176
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_MSB                         183
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_LSB                         176
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_REL_RANGE               183:176
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_REL_MSB                     183
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_REL_LSB                     176
`define DCM_DESKEWTABLEDESC_TLQ0DESKEWCOUNT_RESET_VALUE               8'h93

// macros with short names for field Dcm_DeskewTableDesc.tlq0DeskewCount
`define DCM_DSKWTBLDSC_TLQ0DSKWCNT_RANGE                            183:176
`define DCM_DSKWTBLDSC_TLQ0DSKWCNT_MSB                                  183
`define DCM_DSKWTBLDSC_TLQ0DSKWCNT_LSB                                  176
`define DCM_DSKWTBLDSC_TLQ0DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TLQ0DSKWCNT_RESET_VALUE                        8'h93

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tlq1DeskewCount
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_RANGE                   191:184
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_MSB                         191
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_LSB                         184
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_REL_RANGE               191:184
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_REL_MSB                     191
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_REL_LSB                     184
`define DCM_DESKEWTABLEDESC_TLQ1DESKEWCOUNT_RESET_VALUE               8'h91

// macros with short names for field Dcm_DeskewTableDesc.tlq1DeskewCount
`define DCM_DSKWTBLDSC_TLQ1DSKWCNT_RANGE                            191:184
`define DCM_DSKWTBLDSC_TLQ1DSKWCNT_MSB                                  191
`define DCM_DSKWTBLDSC_TLQ1DSKWCNT_LSB                                  184
`define DCM_DSKWTBLDSC_TLQ1DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TLQ1DSKWCNT_RESET_VALUE                        8'h91

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm9DeskewCount
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_RANGE                   199:192
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_MSB                         199
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_LSB                         192
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_REL_RANGE               199:192
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_REL_MSB                     199
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_REL_LSB                     192
`define DCM_DESKEWTABLEDESC_DMM9DESKEWCOUNT_RESET_VALUE               8'h8f

// macros with short names for field Dcm_DeskewTableDesc.dmm9DeskewCount
`define DCM_DSKWTBLDSC_DMM9DSKWCNT_RANGE                            199:192
`define DCM_DSKWTBLDSC_DMM9DSKWCNT_MSB                                  199
`define DCM_DSKWTBLDSC_DMM9DSKWCNT_LSB                                  192
`define DCM_DSKWTBLDSC_DMM9DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM9DSKWCNT_RESET_VALUE                        8'h8f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fse0DeskewCount
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_RANGE                   207:200
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_MSB                         207
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_LSB                         200
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_REL_RANGE               207:200
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_REL_MSB                     207
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_REL_LSB                     200
`define DCM_DESKEWTABLEDESC_FSE0DESKEWCOUNT_RESET_VALUE               8'h8f

// macros with short names for field Dcm_DeskewTableDesc.fse0DeskewCount
`define DCM_DSKWTBLDSC_FS0DSKWCNT_RANGE                             207:200
`define DCM_DSKWTBLDSC_FS0DSKWCNT_MSB                                   207
`define DCM_DSKWTBLDSC_FS0DSKWCNT_LSB                                   200
`define DCM_DSKWTBLDSC_FS0DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_FS0DSKWCNT_RESET_VALUE                         8'h8f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fse1DeskewCount
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_RANGE                   215:208
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_MSB                         215
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_LSB                         208
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_REL_RANGE               215:208
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_REL_MSB                     215
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_REL_LSB                     208
`define DCM_DESKEWTABLEDESC_FSE1DESKEWCOUNT_RESET_VALUE               8'h8d

// macros with short names for field Dcm_DeskewTableDesc.fse1DeskewCount
`define DCM_DSKWTBLDSC_FS1DSKWCNT_RANGE                             215:208
`define DCM_DSKWTBLDSC_FS1DSKWCNT_MSB                                   215
`define DCM_DSKWTBLDSC_FS1DSKWCNT_LSB                                   208
`define DCM_DSKWTBLDSC_FS1DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_FS1DSKWCNT_RESET_VALUE                         8'h8d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fse2DeskewCount
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_RANGE                   223:216
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_MSB                         223
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_LSB                         216
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_REL_RANGE               223:216
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_REL_MSB                     223
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_REL_LSB                     216
`define DCM_DESKEWTABLEDESC_FSE2DESKEWCOUNT_RESET_VALUE               8'h8d

// macros with short names for field Dcm_DeskewTableDesc.fse2DeskewCount
`define DCM_DSKWTBLDSC_FS2DSKWCNT_RANGE                             223:216
`define DCM_DSKWTBLDSC_FS2DSKWCNT_MSB                                   223
`define DCM_DSKWTBLDSC_FS2DSKWCNT_LSB                                   216
`define DCM_DSKWTBLDSC_FS2DSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_FS2DSKWCNT_RESET_VALUE                         8'h8d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.hsh0DeskewCount
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_RANGE                   231:224
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_MSB                         231
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_LSB                         224
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_REL_RANGE               231:224
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_REL_MSB                     231
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_REL_LSB                     224
`define DCM_DESKEWTABLEDESC_HSH0DESKEWCOUNT_RESET_VALUE               8'h8b

// macros with short names for field Dcm_DeskewTableDesc.hsh0DeskewCount
`define DCM_DSKWTBLDSC_HSH0DSKWCNT_RANGE                            231:224
`define DCM_DSKWTBLDSC_HSH0DSKWCNT_MSB                                  231
`define DCM_DSKWTBLDSC_HSH0DSKWCNT_LSB                                  224
`define DCM_DSKWTBLDSC_HSH0DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_HSH0DSKWCNT_RESET_VALUE                        8'h8b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.hsh1DeskewCount
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_RANGE                   239:232
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_MSB                         239
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_LSB                         232
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_REL_RANGE               239:232
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_REL_MSB                     239
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_REL_LSB                     232
`define DCM_DESKEWTABLEDESC_HSH1DESKEWCOUNT_RESET_VALUE               8'h89

// macros with short names for field Dcm_DeskewTableDesc.hsh1DeskewCount
`define DCM_DSKWTBLDSC_HSH1DSKWCNT_RANGE                            239:232
`define DCM_DSKWTBLDSC_HSH1DSKWCNT_MSB                                  239
`define DCM_DSKWTBLDSC_HSH1DSKWCNT_LSB                                  232
`define DCM_DSKWTBLDSC_HSH1DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_HSH1DSKWCNT_RESET_VALUE                        8'h89

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.hsh2DeskewCount
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_RANGE                   247:240
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_MSB                         247
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_LSB                         240
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_REL_RANGE               247:240
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_REL_MSB                     247
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_REL_LSB                     240
`define DCM_DESKEWTABLEDESC_HSH2DESKEWCOUNT_RESET_VALUE               8'h87

// macros with short names for field Dcm_DeskewTableDesc.hsh2DeskewCount
`define DCM_DSKWTBLDSC_HSH2DSKWCNT_RANGE                            247:240
`define DCM_DSKWTBLDSC_HSH2DSKWCNT_MSB                                  247
`define DCM_DSKWTBLDSC_HSH2DSKWCNT_LSB                                  240
`define DCM_DSKWTBLDSC_HSH2DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_HSH2DSKWCNT_RESET_VALUE                        8'h87

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.hsh3DeskewCount
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_RANGE                   255:248
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_MSB                         255
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_LSB                         248
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_REL_RANGE               255:248
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_REL_MSB                     255
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_REL_LSB                     248
`define DCM_DESKEWTABLEDESC_HSH3DESKEWCOUNT_RESET_VALUE               8'h85

// macros with short names for field Dcm_DeskewTableDesc.hsh3DeskewCount
`define DCM_DSKWTBLDSC_HSH3DSKWCNT_RANGE                            255:248
`define DCM_DSKWTBLDSC_HSH3DSKWCNT_MSB                                  255
`define DCM_DSKWTBLDSC_HSH3DSKWCNT_LSB                                  248
`define DCM_DSKWTBLDSC_HSH3DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_HSH3DSKWCNT_RESET_VALUE                        8'h85

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.hsh4DeskewCount
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_RANGE                   263:256
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_MSB                         263
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_LSB                         256
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_REL_RANGE               263:256
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_REL_MSB                     263
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_REL_LSB                     256
`define DCM_DESKEWTABLEDESC_HSH4DESKEWCOUNT_RESET_VALUE               8'h83

// macros with short names for field Dcm_DeskewTableDesc.hsh4DeskewCount
`define DCM_DSKWTBLDSC_HSH4DSKWCNT_RANGE                            263:256
`define DCM_DSKWTBLDSC_HSH4DSKWCNT_MSB                                  263
`define DCM_DSKWTBLDSC_HSH4DSKWCNT_LSB                                  256
`define DCM_DSKWTBLDSC_HSH4DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_HSH4DSKWCNT_RESET_VALUE                        8'h83

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.oft0DeskewCount
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_RANGE                   271:264
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_MSB                         271
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_LSB                         264
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_REL_RANGE               271:264
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_REL_MSB                     271
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_REL_LSB                     264
`define DCM_DESKEWTABLEDESC_OFT0DESKEWCOUNT_RESET_VALUE               8'h80

// macros with short names for field Dcm_DeskewTableDesc.oft0DeskewCount
`define DCM_DSKWTBLDSC_OFT0DSKWCNT_RANGE                            271:264
`define DCM_DSKWTBLDSC_OFT0DSKWCNT_MSB                                  271
`define DCM_DSKWTBLDSC_OFT0DSKWCNT_LSB                                  264
`define DCM_DSKWTBLDSC_OFT0DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_OFT0DSKWCNT_RESET_VALUE                        8'h80

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.oft1DeskewCount
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_RANGE                   279:272
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_MSB                         279
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_LSB                         272
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_REL_RANGE               279:272
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_REL_MSB                     279
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_REL_LSB                     272
`define DCM_DESKEWTABLEDESC_OFT1DESKEWCOUNT_RESET_VALUE               8'h80

// macros with short names for field Dcm_DeskewTableDesc.oft1DeskewCount
`define DCM_DSKWTBLDSC_OFT1DSKWCNT_RANGE                            279:272
`define DCM_DSKWTBLDSC_OFT1DSKWCNT_MSB                                  279
`define DCM_DSKWTBLDSC_OFT1DSKWCNT_LSB                                  272
`define DCM_DSKWTBLDSC_OFT1DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_OFT1DSKWCNT_RESET_VALUE                        8'h80

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tfq0DeskewCount
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_RANGE                   287:280
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_MSB                         287
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_LSB                         280
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_REL_RANGE               287:280
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_REL_MSB                     287
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_REL_LSB                     280
`define DCM_DESKEWTABLEDESC_TFQ0DESKEWCOUNT_RESET_VALUE               8'h7e

// macros with short names for field Dcm_DeskewTableDesc.tfq0DeskewCount
`define DCM_DSKWTBLDSC_TFQ0DSKWCNT_RANGE                            287:280
`define DCM_DSKWTBLDSC_TFQ0DSKWCNT_MSB                                  287
`define DCM_DSKWTBLDSC_TFQ0DSKWCNT_LSB                                  280
`define DCM_DSKWTBLDSC_TFQ0DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TFQ0DSKWCNT_RESET_VALUE                        8'h7e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.tfq1DeskewCount
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_RANGE                   295:288
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_MSB                         295
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_LSB                         288
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_REL_RANGE               295:288
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_REL_MSB                     295
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_REL_LSB                     288
`define DCM_DESKEWTABLEDESC_TFQ1DESKEWCOUNT_RESET_VALUE               8'h7c

// macros with short names for field Dcm_DeskewTableDesc.tfq1DeskewCount
`define DCM_DSKWTBLDSC_TFQ1DSKWCNT_RANGE                            295:288
`define DCM_DSKWTBLDSC_TFQ1DSKWCNT_MSB                                  295
`define DCM_DSKWTBLDSC_TFQ1DSKWCNT_LSB                                  288
`define DCM_DSKWTBLDSC_TFQ1DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_TFQ1DSKWCNT_RESET_VALUE                        8'h7c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm0DeskewCount
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_RANGE                   303:296
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_MSB                         303
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_LSB                         296
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_REL_RANGE               303:296
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_REL_MSB                     303
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_REL_LSB                     296
`define DCM_DESKEWTABLEDESC_DMM0DESKEWCOUNT_RESET_VALUE               8'h7a

// macros with short names for field Dcm_DeskewTableDesc.dmm0DeskewCount
`define DCM_DSKWTBLDSC_DMM0DSKWCNT_RANGE                            303:296
`define DCM_DSKWTBLDSC_DMM0DSKWCNT_MSB                                  303
`define DCM_DSKWTBLDSC_DMM0DSKWCNT_LSB                                  296
`define DCM_DSKWTBLDSC_DMM0DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM0DSKWCNT_RESET_VALUE                        8'h7a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm1DeskewCount
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_RANGE                   311:304
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_MSB                         311
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_LSB                         304
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_REL_RANGE               311:304
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_REL_MSB                     311
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_REL_LSB                     304
`define DCM_DESKEWTABLEDESC_DMM1DESKEWCOUNT_RESET_VALUE               8'h79

// macros with short names for field Dcm_DeskewTableDesc.dmm1DeskewCount
`define DCM_DSKWTBLDSC_DMM1DSKWCNT_RANGE                            311:304
`define DCM_DSKWTBLDSC_DMM1DSKWCNT_MSB                                  311
`define DCM_DSKWTBLDSC_DMM1DSKWCNT_LSB                                  304
`define DCM_DSKWTBLDSC_DMM1DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM1DSKWCNT_RESET_VALUE                        8'h79

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm2DeskewCount
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_RANGE                   319:312
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_MSB                         319
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_LSB                         312
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_REL_RANGE               319:312
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_REL_MSB                     319
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_REL_LSB                     312
`define DCM_DESKEWTABLEDESC_DMM2DESKEWCOUNT_RESET_VALUE               8'h78

// macros with short names for field Dcm_DeskewTableDesc.dmm2DeskewCount
`define DCM_DSKWTBLDSC_DMM2DSKWCNT_RANGE                            319:312
`define DCM_DSKWTBLDSC_DMM2DSKWCNT_MSB                                  319
`define DCM_DSKWTBLDSC_DMM2DSKWCNT_LSB                                  312
`define DCM_DSKWTBLDSC_DMM2DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM2DSKWCNT_RESET_VALUE                        8'h78

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.pimDeskewCount
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_RANGE                    327:320
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_MSB                          327
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_LSB                          320
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_REL_RANGE                327:320
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_REL_MSB                      327
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_REL_LSB                      320
`define DCM_DESKEWTABLEDESC_PIMDESKEWCOUNT_RESET_VALUE                8'h77

// macros with short names for field Dcm_DeskewTableDesc.pimDeskewCount
`define DCM_DSKWTBLDSC_PMDSKWCNT_RANGE                              327:320
`define DCM_DSKWTBLDSC_PMDSKWCNT_MSB                                    327
`define DCM_DSKWTBLDSC_PMDSKWCNT_LSB                                    320
`define DCM_DSKWTBLDSC_PMDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_PMDSKWCNT_RESET_VALUE                          8'h77

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.supDeskewCount
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_RANGE                    335:328
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_MSB                          335
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_LSB                          328
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_REL_RANGE                335:328
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_REL_MSB                      335
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_REL_LSB                      328
`define DCM_DESKEWTABLEDESC_SUPDESKEWCOUNT_RESET_VALUE                8'h76

// macros with short names for field Dcm_DeskewTableDesc.supDeskewCount
`define DCM_DSKWTBLDSC_SPDSKWCNT_RANGE                              335:328
`define DCM_DSKWTBLDSC_SPDSKWCNT_MSB                                    335
`define DCM_DSKWTBLDSC_SPDSKWCNT_LSB                                    328
`define DCM_DSKWTBLDSC_SPDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_SPDSKWCNT_RESET_VALUE                          8'h76

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm3DeskewCount
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_RANGE                   343:336
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_MSB                         343
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_LSB                         336
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_REL_RANGE               343:336
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_REL_MSB                     343
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_REL_LSB                     336
`define DCM_DESKEWTABLEDESC_DMM3DESKEWCOUNT_RESET_VALUE               8'h73

// macros with short names for field Dcm_DeskewTableDesc.dmm3DeskewCount
`define DCM_DSKWTBLDSC_DMM3DSKWCNT_RANGE                            343:336
`define DCM_DSKWTBLDSC_DMM3DSKWCNT_MSB                                  343
`define DCM_DSKWTBLDSC_DMM3DSKWCNT_LSB                                  336
`define DCM_DSKWTBLDSC_DMM3DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM3DSKWCNT_RESET_VALUE                        8'h73

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm4DeskewCount
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_RANGE                   351:344
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_MSB                         351
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_LSB                         344
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_REL_RANGE               351:344
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_REL_MSB                     351
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_REL_LSB                     344
`define DCM_DESKEWTABLEDESC_DMM4DESKEWCOUNT_RESET_VALUE               8'h72

// macros with short names for field Dcm_DeskewTableDesc.dmm4DeskewCount
`define DCM_DSKWTBLDSC_DMM4DSKWCNT_RANGE                            351:344
`define DCM_DSKWTBLDSC_DMM4DSKWCNT_MSB                                  351
`define DCM_DSKWTBLDSC_DMM4DSKWCNT_LSB                                  344
`define DCM_DSKWTBLDSC_DMM4DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM4DSKWCNT_RESET_VALUE                        8'h72

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm20DeskewCount
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_RANGE                  359:352
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_MSB                        359
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_LSB                        352
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_REL_RANGE              359:352
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_REL_MSB                    359
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_REL_LSB                    352
`define DCM_DESKEWTABLEDESC_DMM20DESKEWCOUNT_RESET_VALUE              8'h71

// macros with short names for field Dcm_DeskewTableDesc.dmm20DeskewCount
`define DCM_DSKWTBLDSC_DMM20DSKWCNT_RANGE                           359:352
`define DCM_DSKWTBLDSC_DMM20DSKWCNT_MSB                                 359
`define DCM_DSKWTBLDSC_DMM20DSKWCNT_LSB                                 352
`define DCM_DSKWTBLDSC_DMM20DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM20DSKWCNT_RESET_VALUE                       8'h71

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm5DeskewCount
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_RANGE                   367:360
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_MSB                         367
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_LSB                         360
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_REL_RANGE               367:360
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_REL_MSB                     367
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_REL_LSB                     360
`define DCM_DESKEWTABLEDESC_DMM5DESKEWCOUNT_RESET_VALUE               8'h70

// macros with short names for field Dcm_DeskewTableDesc.dmm5DeskewCount
`define DCM_DSKWTBLDSC_DMM5DSKWCNT_RANGE                            367:360
`define DCM_DSKWTBLDSC_DMM5DSKWCNT_MSB                                  367
`define DCM_DSKWTBLDSC_DMM5DSKWCNT_LSB                                  360
`define DCM_DSKWTBLDSC_DMM5DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM5DSKWCNT_RESET_VALUE                        8'h70

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.rmuDeskewCount
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_RANGE                    375:368
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_MSB                          375
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_LSB                          368
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_REL_RANGE                375:368
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_REL_MSB                      375
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_REL_LSB                      368
`define DCM_DESKEWTABLEDESC_RMUDESKEWCOUNT_RESET_VALUE                8'h6f

// macros with short names for field Dcm_DeskewTableDesc.rmuDeskewCount
`define DCM_DSKWTBLDSC_RMDSKWCNT_RANGE                              375:368
`define DCM_DSKWTBLDSC_RMDSKWCNT_MSB                                    375
`define DCM_DSKWTBLDSC_RMDSKWCNT_LSB                                    368
`define DCM_DSKWTBLDSC_RMDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_RMDSKWCNT_RESET_VALUE                          8'h6f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.secDeskewCount
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_RANGE                    383:376
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_MSB                          383
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_LSB                          376
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_REL_RANGE                383:376
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_REL_MSB                      383
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_REL_LSB                      376
`define DCM_DESKEWTABLEDESC_SECDESKEWCOUNT_RESET_VALUE                8'h6f

// macros with short names for field Dcm_DeskewTableDesc.secDeskewCount
`define DCM_DSKWTBLDSC_SCDSKWCNT_RANGE                              383:376
`define DCM_DSKWTBLDSC_SCDSKWCNT_MSB                                    383
`define DCM_DSKWTBLDSC_SCDSKWCNT_LSB                                    376
`define DCM_DSKWTBLDSC_SCDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_SCDSKWCNT_RESET_VALUE                          8'h6f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.rreDeskewCount
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_RANGE                    391:384
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_MSB                          391
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_LSB                          384
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_REL_RANGE                391:384
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_REL_MSB                      391
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_REL_LSB                      384
`define DCM_DESKEWTABLEDESC_RREDESKEWCOUNT_RESET_VALUE                8'h6c

// macros with short names for field Dcm_DeskewTableDesc.rreDeskewCount
`define DCM_DSKWTBLDSC_RRDSKWCNT_RANGE                              391:384
`define DCM_DSKWTBLDSC_RRDSKWCNT_MSB                                    391
`define DCM_DSKWTBLDSC_RRDSKWCNT_LSB                                    384
`define DCM_DSKWTBLDSC_RRDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_RRDSKWCNT_RESET_VALUE                          8'h6c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm21DeskewCount
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_RANGE                  399:392
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_MSB                        399
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_LSB                        392
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_REL_RANGE              399:392
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_REL_MSB                    399
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_REL_LSB                    392
`define DCM_DESKEWTABLEDESC_DMM21DESKEWCOUNT_RESET_VALUE              8'h69

// macros with short names for field Dcm_DeskewTableDesc.dmm21DeskewCount
`define DCM_DSKWTBLDSC_DMM21DSKWCNT_RANGE                           399:392
`define DCM_DSKWTBLDSC_DMM21DSKWCNT_MSB                                 399
`define DCM_DSKWTBLDSC_DMM21DSKWCNT_LSB                                 392
`define DCM_DSKWTBLDSC_DMM21DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM21DSKWCNT_RESET_VALUE                       8'h69

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.nifDeskewCount
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_RANGE                    407:400
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_MSB                          407
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_LSB                          400
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_REL_RANGE                407:400
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_REL_MSB                      407
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_REL_LSB                      400
`define DCM_DESKEWTABLEDESC_NIFDESKEWCOUNT_RESET_VALUE                8'h6a

// macros with short names for field Dcm_DeskewTableDesc.nifDeskewCount
`define DCM_DSKWTBLDSC_NFDSKWCNT_RANGE                              407:400
`define DCM_DSKWTBLDSC_NFDSKWCNT_MSB                                    407
`define DCM_DSKWTBLDSC_NFDSKWCNT_LSB                                    400
`define DCM_DSKWTBLDSC_NFDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_NFDSKWCNT_RESET_VALUE                          8'h6a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ipfDeskewCount
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_RANGE                    415:408
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_MSB                          415
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_LSB                          408
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_REL_RANGE                415:408
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_REL_MSB                      415
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_REL_LSB                      408
`define DCM_DESKEWTABLEDESC_IPFDESKEWCOUNT_RESET_VALUE                8'h66

// macros with short names for field Dcm_DeskewTableDesc.ipfDeskewCount
`define DCM_DSKWTBLDSC_IPFDSKWCNT_RANGE                             415:408
`define DCM_DSKWTBLDSC_IPFDSKWCNT_MSB                                   415
`define DCM_DSKWTBLDSC_IPFDSKWCNT_LSB                                   408
`define DCM_DSKWTBLDSC_IPFDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_IPFDSKWCNT_RESET_VALUE                         8'h66

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm23DeskewCount
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_RANGE                  423:416
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_MSB                        423
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_LSB                        416
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_REL_RANGE              423:416
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_REL_MSB                    423
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_REL_LSB                    416
`define DCM_DESKEWTABLEDESC_DMM23DESKEWCOUNT_RESET_VALUE              8'h64

// macros with short names for field Dcm_DeskewTableDesc.dmm23DeskewCount
`define DCM_DSKWTBLDSC_DMM23DSKWCNT_RANGE                           423:416
`define DCM_DSKWTBLDSC_DMM23DSKWCNT_MSB                                 423
`define DCM_DSKWTBLDSC_DMM23DSKWCNT_LSB                                 416
`define DCM_DSKWTBLDSC_DMM23DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM23DSKWCNT_RESET_VALUE                       8'h64

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.mscIngressDeskewCount
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_RANGE             431:424
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_MSB                   431
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_LSB                   424
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_WIDTH                   8
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_REL_RANGE         431:424
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_REL_MSB               431
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_REL_LSB               424
`define DCM_DESKEWTABLEDESC_MSCINGRESSDESKEWCOUNT_RESET_VALUE         8'h63

// macros with short names for field Dcm_DeskewTableDesc.mscIngressDeskewCount
`define DCM_DSKWTBLDSC_MSCINGRDSKWCNT_RANGE                         431:424
`define DCM_DSKWTBLDSC_MSCINGRDSKWCNT_MSB                               431
`define DCM_DSKWTBLDSC_MSCINGRDSKWCNT_LSB                               424
`define DCM_DSKWTBLDSC_MSCINGRDSKWCNT_WIDTH                               8
`define DCM_DSKWTBLDSC_MSCINGRDSKWCNT_RESET_VALUE                     8'h63

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm24DeskewCount
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_RANGE                  439:432
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_MSB                        439
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_LSB                        432
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_REL_RANGE              439:432
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_REL_MSB                    439
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_REL_LSB                    432
`define DCM_DESKEWTABLEDESC_DMM24DESKEWCOUNT_RESET_VALUE              8'h61

// macros with short names for field Dcm_DeskewTableDesc.dmm24DeskewCount
`define DCM_DSKWTBLDSC_DMM24DSKWCNT_RANGE                           439:432
`define DCM_DSKWTBLDSC_DMM24DSKWCNT_MSB                                 439
`define DCM_DSKWTBLDSC_DMM24DSKWCNT_LSB                                 432
`define DCM_DSKWTBLDSC_DMM24DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM24DSKWCNT_RESET_VALUE                       8'h61

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fpeIngressDeskewCount
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_RANGE             447:440
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_MSB                   447
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_LSB                   440
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_WIDTH                   8
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_REL_RANGE         447:440
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_REL_MSB               447
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_REL_LSB               440
`define DCM_DESKEWTABLEDESC_FPEINGRESSDESKEWCOUNT_RESET_VALUE         8'h62

// macros with short names for field Dcm_DeskewTableDesc.fpeIngressDeskewCount
`define DCM_DSKWTBLDSC_FPINGRDSKWCNT_RANGE                          447:440
`define DCM_DSKWTBLDSC_FPINGRDSKWCNT_MSB                                447
`define DCM_DSKWTBLDSC_FPINGRDSKWCNT_LSB                                440
`define DCM_DSKWTBLDSC_FPINGRDSKWCNT_WIDTH                                8
`define DCM_DSKWTBLDSC_FPINGRDSKWCNT_RESET_VALUE                      8'h62

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.cmmDeskewCount
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_RANGE                    455:448
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_MSB                          455
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_LSB                          448
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_REL_RANGE                455:448
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_REL_MSB                      455
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_REL_LSB                      448
`define DCM_DESKEWTABLEDESC_CMMDESKEWCOUNT_RESET_VALUE                8'h60

// macros with short names for field Dcm_DeskewTableDesc.cmmDeskewCount
`define DCM_DSKWTBLDSC_CMMDSKWCNT_RANGE                             455:448
`define DCM_DSKWTBLDSC_CMMDSKWCNT_MSB                                   455
`define DCM_DSKWTBLDSC_CMMDSKWCNT_LSB                                   448
`define DCM_DSKWTBLDSC_CMMDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_CMMDSKWCNT_RESET_VALUE                         8'h60

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm19DeskewCount
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_RANGE                  463:456
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_MSB                        463
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_LSB                        456
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_REL_RANGE              463:456
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_REL_MSB                    463
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_REL_LSB                    456
`define DCM_DESKEWTABLEDESC_DMM19DESKEWCOUNT_RESET_VALUE              8'h5c

// macros with short names for field Dcm_DeskewTableDesc.dmm19DeskewCount
`define DCM_DSKWTBLDSC_DMM19DSKWCNT_RANGE                           463:456
`define DCM_DSKWTBLDSC_DMM19DSKWCNT_MSB                                 463
`define DCM_DSKWTBLDSC_DMM19DSKWCNT_LSB                                 456
`define DCM_DSKWTBLDSC_DMM19DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM19DSKWCNT_RESET_VALUE                       8'h5c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ippDeskewCount
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_RANGE                    471:464
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_MSB                          471
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_LSB                          464
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_REL_RANGE                471:464
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_REL_MSB                      471
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_REL_LSB                      464
`define DCM_DESKEWTABLEDESC_IPPDESKEWCOUNT_RESET_VALUE                8'h5d

// macros with short names for field Dcm_DeskewTableDesc.ippDeskewCount
`define DCM_DSKWTBLDSC_IPPDSKWCNT_RANGE                             471:464
`define DCM_DSKWTBLDSC_IPPDSKWCNT_MSB                                   471
`define DCM_DSKWTBLDSC_IPPDSKWCNT_LSB                                   464
`define DCM_DSKWTBLDSC_IPPDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_IPPDSKWCNT_RESET_VALUE                         8'h5d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm18DeskewCount
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_RANGE                  479:472
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_MSB                        479
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_LSB                        472
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_REL_RANGE              479:472
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_REL_MSB                    479
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_REL_LSB                    472
`define DCM_DESKEWTABLEDESC_DMM18DESKEWCOUNT_RESET_VALUE              8'h59

// macros with short names for field Dcm_DeskewTableDesc.dmm18DeskewCount
`define DCM_DSKWTBLDSC_DMM18DSKWCNT_RANGE                           479:472
`define DCM_DSKWTBLDSC_DMM18DSKWCNT_MSB                                 479
`define DCM_DSKWTBLDSC_DMM18DSKWCNT_LSB                                 472
`define DCM_DSKWTBLDSC_DMM18DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM18DSKWCNT_RESET_VALUE                       8'h59

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps0DeskewCount
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_RANGE                   487:480
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_MSB                         487
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_LSB                         480
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_REL_RANGE               487:480
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_REL_MSB                     487
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_REL_LSB                     480
`define DCM_DESKEWTABLEDESC_FPS0DESKEWCOUNT_RESET_VALUE               8'h59

// macros with short names for field Dcm_DeskewTableDesc.fps0DeskewCount
`define DCM_DSKWTBLDSC_FPS0DSKWCNT_RANGE                            487:480
`define DCM_DSKWTBLDSC_FPS0DSKWCNT_MSB                                  487
`define DCM_DSKWTBLDSC_FPS0DSKWCNT_LSB                                  480
`define DCM_DSKWTBLDSC_FPS0DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS0DSKWCNT_RESET_VALUE                        8'h59

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.ileDeskewCount
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_RANGE                    495:488
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_MSB                          495
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_LSB                          488
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_REL_RANGE                495:488
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_REL_MSB                      495
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_REL_LSB                      488
`define DCM_DESKEWTABLEDESC_ILEDESKEWCOUNT_RESET_VALUE                8'h58

// macros with short names for field Dcm_DeskewTableDesc.ileDeskewCount
`define DCM_DSKWTBLDSC_ILDSKWCNT_RANGE                              495:488
`define DCM_DSKWTBLDSC_ILDSKWCNT_MSB                                    495
`define DCM_DSKWTBLDSC_ILDSKWCNT_LSB                                    488
`define DCM_DSKWTBLDSC_ILDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_ILDSKWCNT_RESET_VALUE                          8'h58

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps1DeskewCount
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_RANGE                   503:496
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_MSB                         503
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_LSB                         496
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_REL_RANGE               503:496
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_REL_MSB                     503
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_REL_LSB                     496
`define DCM_DESKEWTABLEDESC_FPS1DESKEWCOUNT_RESET_VALUE               8'h55

// macros with short names for field Dcm_DeskewTableDesc.fps1DeskewCount
`define DCM_DSKWTBLDSC_FPS1DSKWCNT_RANGE                            503:496
`define DCM_DSKWTBLDSC_FPS1DSKWCNT_MSB                                  503
`define DCM_DSKWTBLDSC_FPS1DSKWCNT_LSB                                  496
`define DCM_DSKWTBLDSC_FPS1DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS1DSKWCNT_RESET_VALUE                        8'h55

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps2DeskewCount
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_RANGE                   511:504
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_MSB                         511
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_LSB                         504
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_REL_RANGE               511:504
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_REL_MSB                     511
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_REL_LSB                     504
`define DCM_DESKEWTABLEDESC_FPS2DESKEWCOUNT_RESET_VALUE               8'h53

// macros with short names for field Dcm_DeskewTableDesc.fps2DeskewCount
`define DCM_DSKWTBLDSC_FPS2DSKWCNT_RANGE                            511:504
`define DCM_DSKWTBLDSC_FPS2DSKWCNT_MSB                                  511
`define DCM_DSKWTBLDSC_FPS2DSKWCNT_LSB                                  504
`define DCM_DSKWTBLDSC_FPS2DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS2DSKWCNT_RESET_VALUE                        8'h53

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps3DeskewCount
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_RANGE                   519:512
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_MSB                         519
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_LSB                         512
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_REL_RANGE               519:512
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_REL_MSB                     519
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_REL_LSB                     512
`define DCM_DESKEWTABLEDESC_FPS3DESKEWCOUNT_RESET_VALUE               8'h51

// macros with short names for field Dcm_DeskewTableDesc.fps3DeskewCount
`define DCM_DSKWTBLDSC_FPS3DSKWCNT_RANGE                            519:512
`define DCM_DSKWTBLDSC_FPS3DSKWCNT_MSB                                  519
`define DCM_DSKWTBLDSC_FPS3DSKWCNT_LSB                                  512
`define DCM_DSKWTBLDSC_FPS3DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS3DSKWCNT_RESET_VALUE                        8'h51

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps4DeskewCount
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_RANGE                   527:520
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_MSB                         527
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_LSB                         520
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_REL_RANGE               527:520
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_REL_MSB                     527
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_REL_LSB                     520
`define DCM_DESKEWTABLEDESC_FPS4DESKEWCOUNT_RESET_VALUE               8'h4f

// macros with short names for field Dcm_DeskewTableDesc.fps4DeskewCount
`define DCM_DSKWTBLDSC_FPS4DSKWCNT_RANGE                            527:520
`define DCM_DSKWTBLDSC_FPS4DSKWCNT_MSB                                  527
`define DCM_DSKWTBLDSC_FPS4DSKWCNT_LSB                                  520
`define DCM_DSKWTBLDSC_FPS4DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS4DSKWCNT_RESET_VALUE                        8'h4f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps5DeskewCount
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_RANGE                   535:528
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_MSB                         535
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_LSB                         528
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_REL_RANGE               535:528
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_REL_MSB                     535
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_REL_LSB                     528
`define DCM_DESKEWTABLEDESC_FPS5DESKEWCOUNT_RESET_VALUE               8'h4d

// macros with short names for field Dcm_DeskewTableDesc.fps5DeskewCount
`define DCM_DSKWTBLDSC_FPS5DSKWCNT_RANGE                            535:528
`define DCM_DSKWTBLDSC_FPS5DSKWCNT_MSB                                  535
`define DCM_DSKWTBLDSC_FPS5DSKWCNT_LSB                                  528
`define DCM_DSKWTBLDSC_FPS5DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS5DSKWCNT_RESET_VALUE                        8'h4d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps6DeskewCount
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_RANGE                   543:536
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_MSB                         543
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_LSB                         536
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_REL_RANGE               543:536
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_REL_MSB                     543
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_REL_LSB                     536
`define DCM_DESKEWTABLEDESC_FPS6DESKEWCOUNT_RESET_VALUE               8'h4b

// macros with short names for field Dcm_DeskewTableDesc.fps6DeskewCount
`define DCM_DSKWTBLDSC_FPS6DSKWCNT_RANGE                            543:536
`define DCM_DSKWTBLDSC_FPS6DSKWCNT_MSB                                  543
`define DCM_DSKWTBLDSC_FPS6DSKWCNT_LSB                                  536
`define DCM_DSKWTBLDSC_FPS6DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS6DSKWCNT_RESET_VALUE                        8'h4b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps7DeskewCount
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_RANGE                   551:544
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_MSB                         551
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_LSB                         544
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_REL_RANGE               551:544
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_REL_MSB                     551
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_REL_LSB                     544
`define DCM_DESKEWTABLEDESC_FPS7DESKEWCOUNT_RESET_VALUE               8'h49

// macros with short names for field Dcm_DeskewTableDesc.fps7DeskewCount
`define DCM_DSKWTBLDSC_FPS7DSKWCNT_RANGE                            551:544
`define DCM_DSKWTBLDSC_FPS7DSKWCNT_MSB                                  551
`define DCM_DSKWTBLDSC_FPS7DSKWCNT_LSB                                  544
`define DCM_DSKWTBLDSC_FPS7DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS7DSKWCNT_RESET_VALUE                        8'h49

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps8DeskewCount
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_RANGE                   559:552
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_MSB                         559
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_LSB                         552
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_REL_RANGE               559:552
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_REL_MSB                     559
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_REL_LSB                     552
`define DCM_DESKEWTABLEDESC_FPS8DESKEWCOUNT_RESET_VALUE               8'h47

// macros with short names for field Dcm_DeskewTableDesc.fps8DeskewCount
`define DCM_DSKWTBLDSC_FPS8DSKWCNT_RANGE                            559:552
`define DCM_DSKWTBLDSC_FPS8DSKWCNT_MSB                                  559
`define DCM_DSKWTBLDSC_FPS8DSKWCNT_LSB                                  552
`define DCM_DSKWTBLDSC_FPS8DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS8DSKWCNT_RESET_VALUE                        8'h47

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps9DeskewCount
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_RANGE                   567:560
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_MSB                         567
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_LSB                         560
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_REL_RANGE               567:560
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_REL_MSB                     567
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_REL_LSB                     560
`define DCM_DESKEWTABLEDESC_FPS9DESKEWCOUNT_RESET_VALUE               8'h45

// macros with short names for field Dcm_DeskewTableDesc.fps9DeskewCount
`define DCM_DSKWTBLDSC_FPS9DSKWCNT_RANGE                            567:560
`define DCM_DSKWTBLDSC_FPS9DSKWCNT_MSB                                  567
`define DCM_DSKWTBLDSC_FPS9DSKWCNT_LSB                                  560
`define DCM_DSKWTBLDSC_FPS9DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_FPS9DSKWCNT_RESET_VALUE                        8'h45

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps10DeskewCount
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_RANGE                  575:568
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_MSB                        575
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_LSB                        568
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_REL_RANGE              575:568
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_REL_MSB                    575
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_REL_LSB                    568
`define DCM_DESKEWTABLEDESC_FPS10DESKEWCOUNT_RESET_VALUE              8'h43

// macros with short names for field Dcm_DeskewTableDesc.fps10DeskewCount
`define DCM_DSKWTBLDSC_FPS10DSKWCNT_RANGE                           575:568
`define DCM_DSKWTBLDSC_FPS10DSKWCNT_MSB                                 575
`define DCM_DSKWTBLDSC_FPS10DSKWCNT_LSB                                 568
`define DCM_DSKWTBLDSC_FPS10DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS10DSKWCNT_RESET_VALUE                       8'h43

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps11DeskewCount
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_RANGE                  583:576
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_MSB                        583
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_LSB                        576
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_REL_RANGE              583:576
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_REL_MSB                    583
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_REL_LSB                    576
`define DCM_DESKEWTABLEDESC_FPS11DESKEWCOUNT_RESET_VALUE              8'h41

// macros with short names for field Dcm_DeskewTableDesc.fps11DeskewCount
`define DCM_DSKWTBLDSC_FPS11DSKWCNT_RANGE                           583:576
`define DCM_DSKWTBLDSC_FPS11DSKWCNT_MSB                                 583
`define DCM_DSKWTBLDSC_FPS11DSKWCNT_LSB                                 576
`define DCM_DSKWTBLDSC_FPS11DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS11DSKWCNT_RESET_VALUE                       8'h41

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps12DeskewCount
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_RANGE                  591:584
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_MSB                        591
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_LSB                        584
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_REL_RANGE              591:584
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_REL_MSB                    591
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_REL_LSB                    584
`define DCM_DESKEWTABLEDESC_FPS12DESKEWCOUNT_RESET_VALUE              8'h3f

// macros with short names for field Dcm_DeskewTableDesc.fps12DeskewCount
`define DCM_DSKWTBLDSC_FPS12DSKWCNT_RANGE                           591:584
`define DCM_DSKWTBLDSC_FPS12DSKWCNT_MSB                                 591
`define DCM_DSKWTBLDSC_FPS12DSKWCNT_LSB                                 584
`define DCM_DSKWTBLDSC_FPS12DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS12DSKWCNT_RESET_VALUE                       8'h3f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps13DeskewCount
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_RANGE                  599:592
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_MSB                        599
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_LSB                        592
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_REL_RANGE              599:592
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_REL_MSB                    599
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_REL_LSB                    592
`define DCM_DESKEWTABLEDESC_FPS13DESKEWCOUNT_RESET_VALUE              8'h3d

// macros with short names for field Dcm_DeskewTableDesc.fps13DeskewCount
`define DCM_DSKWTBLDSC_FPS13DSKWCNT_RANGE                           599:592
`define DCM_DSKWTBLDSC_FPS13DSKWCNT_MSB                                 599
`define DCM_DSKWTBLDSC_FPS13DSKWCNT_LSB                                 592
`define DCM_DSKWTBLDSC_FPS13DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS13DSKWCNT_RESET_VALUE                       8'h3d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps14DeskewCount
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_RANGE                  607:600
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_MSB                        607
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_LSB                        600
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_REL_RANGE              607:600
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_REL_MSB                    607
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_REL_LSB                    600
`define DCM_DESKEWTABLEDESC_FPS14DESKEWCOUNT_RESET_VALUE              8'h3b

// macros with short names for field Dcm_DeskewTableDesc.fps14DeskewCount
`define DCM_DSKWTBLDSC_FPS14DSKWCNT_RANGE                           607:600
`define DCM_DSKWTBLDSC_FPS14DSKWCNT_MSB                                 607
`define DCM_DSKWTBLDSC_FPS14DSKWCNT_LSB                                 600
`define DCM_DSKWTBLDSC_FPS14DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS14DSKWCNT_RESET_VALUE                       8'h3b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.igrDeskewCount
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_RANGE                    615:608
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_MSB                          615
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_LSB                          608
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_REL_RANGE                615:608
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_REL_MSB                      615
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_REL_LSB                      608
`define DCM_DESKEWTABLEDESC_IGRDESKEWCOUNT_RESET_VALUE                8'h3a

// macros with short names for field Dcm_DeskewTableDesc.igrDeskewCount
`define DCM_DSKWTBLDSC_IGRDSKWCNT_RANGE                             615:608
`define DCM_DSKWTBLDSC_IGRDSKWCNT_MSB                                   615
`define DCM_DSKWTBLDSC_IGRDSKWCNT_LSB                                   608
`define DCM_DSKWTBLDSC_IGRDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_IGRDSKWCNT_RESET_VALUE                         8'h3a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm10DeskewCount
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_RANGE                  623:616
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_MSB                        623
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_LSB                        616
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_REL_RANGE              623:616
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_REL_MSB                    623
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_REL_LSB                    616
`define DCM_DESKEWTABLEDESC_DMM10DESKEWCOUNT_RESET_VALUE              8'h36

// macros with short names for field Dcm_DeskewTableDesc.dmm10DeskewCount
`define DCM_DSKWTBLDSC_DMM10DSKWCNT_RANGE                           623:616
`define DCM_DSKWTBLDSC_DMM10DSKWCNT_MSB                                 623
`define DCM_DSKWTBLDSC_DMM10DSKWCNT_LSB                                 616
`define DCM_DSKWTBLDSC_DMM10DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM10DSKWCNT_RESET_VALUE                       8'h36

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.iqsDeskewCount
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_RANGE                    631:624
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_MSB                          631
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_LSB                          624
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_REL_RANGE                631:624
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_REL_MSB                      631
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_REL_LSB                      624
`define DCM_DESKEWTABLEDESC_IQSDESKEWCOUNT_RESET_VALUE                8'h35

// macros with short names for field Dcm_DeskewTableDesc.iqsDeskewCount
`define DCM_DSKWTBLDSC_IQSDSKWCNT_RANGE                             631:624
`define DCM_DSKWTBLDSC_IQSDSKWCNT_MSB                                   631
`define DCM_DSKWTBLDSC_IQSDSKWCNT_LSB                                   624
`define DCM_DSKWTBLDSC_IQSDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_IQSDSKWCNT_RESET_VALUE                         8'h35

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.sqsDeskewCount
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_RANGE                    639:632
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_MSB                          639
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_LSB                          632
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_REL_RANGE                639:632
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_REL_MSB                      639
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_REL_LSB                      632
`define DCM_DESKEWTABLEDESC_SQSDESKEWCOUNT_RESET_VALUE                8'h33

// macros with short names for field Dcm_DeskewTableDesc.sqsDeskewCount
`define DCM_DSKWTBLDSC_SQSDSKWCNT_RANGE                             639:632
`define DCM_DSKWTBLDSC_SQSDSKWCNT_MSB                                   639
`define DCM_DSKWTBLDSC_SQSDSKWCNT_LSB                                   632
`define DCM_DSKWTBLDSC_SQSDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_SQSDSKWCNT_RESET_VALUE                         8'h33

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.aqmDeskewCount
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_RANGE                    647:640
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_MSB                          647
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_LSB                          640
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_REL_RANGE                647:640
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_REL_MSB                      647
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_REL_LSB                      640
`define DCM_DESKEWTABLEDESC_AQMDESKEWCOUNT_RESET_VALUE                8'h33

// macros with short names for field Dcm_DeskewTableDesc.aqmDeskewCount
`define DCM_DSKWTBLDSC_AQMDSKWCNT_RANGE                             647:640
`define DCM_DSKWTBLDSC_AQMDSKWCNT_MSB                                   647
`define DCM_DSKWTBLDSC_AQMDSKWCNT_LSB                                   640
`define DCM_DSKWTBLDSC_AQMDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_AQMDSKWCNT_RESET_VALUE                         8'h33

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.eqcDeskewCount
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_RANGE                    655:648
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_MSB                          655
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_LSB                          648
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_REL_RANGE                655:648
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_REL_MSB                      655
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_REL_LSB                      648
`define DCM_DESKEWTABLEDESC_EQCDESKEWCOUNT_RESET_VALUE                8'h2f

// macros with short names for field Dcm_DeskewTableDesc.eqcDeskewCount
`define DCM_DSKWTBLDSC_EQCDSKWCNT_RANGE                             655:648
`define DCM_DSKWTBLDSC_EQCDSKWCNT_MSB                                   655
`define DCM_DSKWTBLDSC_EQCDSKWCNT_LSB                                   648
`define DCM_DSKWTBLDSC_EQCDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_EQCDSKWCNT_RESET_VALUE                         8'h2f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.esmDeskewCount
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_RANGE                    663:656
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_MSB                          663
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_LSB                          656
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_REL_RANGE                663:656
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_REL_MSB                      663
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_REL_LSB                      656
`define DCM_DESKEWTABLEDESC_ESMDESKEWCOUNT_RESET_VALUE                8'h2d

// macros with short names for field Dcm_DeskewTableDesc.esmDeskewCount
`define DCM_DSKWTBLDSC_ESMDSKWCNT_RANGE                             663:656
`define DCM_DSKWTBLDSC_ESMDSKWCNT_MSB                                   663
`define DCM_DSKWTBLDSC_ESMDSKWCNT_LSB                                   656
`define DCM_DSKWTBLDSC_ESMDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_ESMDSKWCNT_RESET_VALUE                         8'h2d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.pbcDeskewCount
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_RANGE                    671:664
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_MSB                          671
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_LSB                          664
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_REL_RANGE                671:664
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_REL_MSB                      671
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_REL_LSB                      664
`define DCM_DESKEWTABLEDESC_PBCDESKEWCOUNT_RESET_VALUE                8'h2d

// macros with short names for field Dcm_DeskewTableDesc.pbcDeskewCount
`define DCM_DSKWTBLDSC_PBCDSKWCNT_RANGE                             671:664
`define DCM_DSKWTBLDSC_PBCDSKWCNT_MSB                                   671
`define DCM_DSKWTBLDSC_PBCDSKWCNT_LSB                                   664
`define DCM_DSKWTBLDSC_PBCDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_PBCDSKWCNT_RESET_VALUE                         8'h2d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm15DeskewCount
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_RANGE                  679:672
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_MSB                        679
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_LSB                        672
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_REL_RANGE              679:672
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_REL_MSB                    679
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_REL_LSB                    672
`define DCM_DESKEWTABLEDESC_DMM15DESKEWCOUNT_RESET_VALUE              8'h29

// macros with short names for field Dcm_DeskewTableDesc.dmm15DeskewCount
`define DCM_DSKWTBLDSC_DMM15DSKWCNT_RANGE                           679:672
`define DCM_DSKWTBLDSC_DMM15DSKWCNT_MSB                                 679
`define DCM_DSKWTBLDSC_DMM15DSKWCNT_LSB                                 672
`define DCM_DSKWTBLDSC_DMM15DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM15DSKWCNT_RESET_VALUE                       8'h29

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.sifDeskewCount
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_RANGE                    687:680
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_MSB                          687
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_LSB                          680
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_REL_RANGE                687:680
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_REL_MSB                      687
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_REL_LSB                      680
`define DCM_DESKEWTABLEDESC_SIFDESKEWCOUNT_RESET_VALUE                8'h2a

// macros with short names for field Dcm_DeskewTableDesc.sifDeskewCount
`define DCM_DSKWTBLDSC_SFDSKWCNT_RANGE                              687:680
`define DCM_DSKWTBLDSC_SFDSKWCNT_MSB                                    687
`define DCM_DSKWTBLDSC_SFDSKWCNT_LSB                                    680
`define DCM_DSKWTBLDSC_SFDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_SFDSKWCNT_RESET_VALUE                          8'h2a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm22DeskewCount
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_RANGE                  695:688
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_MSB                        695
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_LSB                        688
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_REL_RANGE              695:688
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_REL_MSB                    695
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_REL_LSB                    688
`define DCM_DESKEWTABLEDESC_DMM22DESKEWCOUNT_RESET_VALUE              8'h25

// macros with short names for field Dcm_DeskewTableDesc.dmm22DeskewCount
`define DCM_DSKWTBLDSC_DMM22DSKWCNT_RANGE                           695:688
`define DCM_DSKWTBLDSC_DMM22DSKWCNT_MSB                                 695
`define DCM_DSKWTBLDSC_DMM22DSKWCNT_LSB                                 688
`define DCM_DSKWTBLDSC_DMM22DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM22DSKWCNT_RESET_VALUE                       8'h25

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm8DeskewCount
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_RANGE                   703:696
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_MSB                         703
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_LSB                         696
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_REL_RANGE               703:696
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_REL_MSB                     703
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_REL_LSB                     696
`define DCM_DESKEWTABLEDESC_DMM8DESKEWCOUNT_RESET_VALUE               8'h24

// macros with short names for field Dcm_DeskewTableDesc.dmm8DeskewCount
`define DCM_DSKWTBLDSC_DMM8DSKWCNT_RANGE                            703:696
`define DCM_DSKWTBLDSC_DMM8DSKWCNT_MSB                                  703
`define DCM_DSKWTBLDSC_DMM8DSKWCNT_LSB                                  696
`define DCM_DSKWTBLDSC_DMM8DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM8DSKWCNT_RESET_VALUE                        8'h24

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fpeEgressDeskewCount
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_RANGE              711:704
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_MSB                    711
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_LSB                    704
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_WIDTH                    8
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_REL_RANGE          711:704
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_REL_MSB                711
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_REL_LSB                704
`define DCM_DESKEWTABLEDESC_FPEEGRESSDESKEWCOUNT_RESET_VALUE          8'h25

// macros with short names for field Dcm_DeskewTableDesc.fpeEgressDeskewCount
`define DCM_DSKWTBLDSC_FPEGRSDSKWCNT_RANGE                          711:704
`define DCM_DSKWTBLDSC_FPEGRSDSKWCNT_MSB                                711
`define DCM_DSKWTBLDSC_FPEGRSDSKWCNT_LSB                                704
`define DCM_DSKWTBLDSC_FPEGRSDSKWCNT_WIDTH                                8
`define DCM_DSKWTBLDSC_FPEGRSDSKWCNT_RESET_VALUE                      8'h25

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm25DeskewCount
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_RANGE                  719:712
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_MSB                        719
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_LSB                        712
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_REL_RANGE              719:712
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_REL_MSB                    719
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_REL_LSB                    712
`define DCM_DESKEWTABLEDESC_DMM25DESKEWCOUNT_RESET_VALUE              8'h21

// macros with short names for field Dcm_DeskewTableDesc.dmm25DeskewCount
`define DCM_DSKWTBLDSC_DMM25DSKWCNT_RANGE                           719:712
`define DCM_DSKWTBLDSC_DMM25DSKWCNT_MSB                                 719
`define DCM_DSKWTBLDSC_DMM25DSKWCNT_LSB                                 712
`define DCM_DSKWTBLDSC_DMM25DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM25DSKWCNT_RESET_VALUE                       8'h21

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm14DeskewCount
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_RANGE                  727:720
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_MSB                        727
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_LSB                        720
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_REL_RANGE              727:720
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_REL_MSB                    727
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_REL_LSB                    720
`define DCM_DESKEWTABLEDESC_DMM14DESKEWCOUNT_RESET_VALUE              8'h20

// macros with short names for field Dcm_DeskewTableDesc.dmm14DeskewCount
`define DCM_DSKWTBLDSC_DMM14DSKWCNT_RANGE                           727:720
`define DCM_DSKWTBLDSC_DMM14DSKWCNT_MSB                                 727
`define DCM_DSKWTBLDSC_DMM14DSKWCNT_LSB                                 720
`define DCM_DSKWTBLDSC_DMM14DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM14DSKWCNT_RESET_VALUE                       8'h20

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.frwDeskewCount
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_RANGE                    735:728
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_MSB                          735
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_LSB                          728
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_REL_RANGE                735:728
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_REL_MSB                      735
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_REL_LSB                      728
`define DCM_DESKEWTABLEDESC_FRWDESKEWCOUNT_RESET_VALUE                8'h21

// macros with short names for field Dcm_DeskewTableDesc.frwDeskewCount
`define DCM_DSKWTBLDSC_FRWDSKWCNT_RANGE                             735:728
`define DCM_DSKWTBLDSC_FRWDSKWCNT_MSB                                   735
`define DCM_DSKWTBLDSC_FRWDSKWCNT_LSB                                   728
`define DCM_DSKWTBLDSC_FRWDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_FRWDSKWCNT_RESET_VALUE                         8'h21

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm16DeskewCount
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_RANGE                  743:736
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_MSB                        743
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_LSB                        736
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_REL_RANGE              743:736
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_REL_MSB                    743
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_REL_LSB                    736
`define DCM_DESKEWTABLEDESC_DMM16DESKEWCOUNT_RESET_VALUE              8'h1d

// macros with short names for field Dcm_DeskewTableDesc.dmm16DeskewCount
`define DCM_DSKWTBLDSC_DMM16DSKWCNT_RANGE                           743:736
`define DCM_DSKWTBLDSC_DMM16DSKWCNT_MSB                                 743
`define DCM_DSKWTBLDSC_DMM16DSKWCNT_LSB                                 736
`define DCM_DSKWTBLDSC_DMM16DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM16DSKWCNT_RESET_VALUE                       8'h1d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.eppDeskewCount
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_RANGE                    751:744
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_MSB                          751
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_LSB                          744
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_REL_RANGE                751:744
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_REL_MSB                      751
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_REL_LSB                      744
`define DCM_DESKEWTABLEDESC_EPPDESKEWCOUNT_RESET_VALUE                8'h1e

// macros with short names for field Dcm_DeskewTableDesc.eppDeskewCount
`define DCM_DSKWTBLDSC_EPPDSKWCNT_RANGE                             751:744
`define DCM_DSKWTBLDSC_EPPDSKWCNT_MSB                                   751
`define DCM_DSKWTBLDSC_EPPDSKWCNT_LSB                                   744
`define DCM_DSKWTBLDSC_EPPDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_EPPDSKWCNT_RESET_VALUE                         8'h1e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps15DeskewCount
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_RANGE                  759:752
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_MSB                        759
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_LSB                        752
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_REL_RANGE              759:752
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_REL_MSB                    759
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_REL_LSB                    752
`define DCM_DESKEWTABLEDESC_FPS15DESKEWCOUNT_RESET_VALUE              8'h1b

// macros with short names for field Dcm_DeskewTableDesc.fps15DeskewCount
`define DCM_DSKWTBLDSC_FPS15DSKWCNT_RANGE                           759:752
`define DCM_DSKWTBLDSC_FPS15DSKWCNT_MSB                                 759
`define DCM_DSKWTBLDSC_FPS15DSKWCNT_LSB                                 752
`define DCM_DSKWTBLDSC_FPS15DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS15DSKWCNT_RESET_VALUE                       8'h1b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.eleDeskewCount
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_RANGE                    767:760
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_MSB                          767
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_LSB                          760
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_REL_RANGE                767:760
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_REL_MSB                      767
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_REL_LSB                      760
`define DCM_DESKEWTABLEDESC_ELEDESKEWCOUNT_RESET_VALUE                8'h1a

// macros with short names for field Dcm_DeskewTableDesc.eleDeskewCount
`define DCM_DSKWTBLDSC_ELDSKWCNT_RANGE                              767:760
`define DCM_DSKWTBLDSC_ELDSKWCNT_MSB                                    767
`define DCM_DSKWTBLDSC_ELDSKWCNT_LSB                                    760
`define DCM_DSKWTBLDSC_ELDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_ELDSKWCNT_RESET_VALUE                          8'h1a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps16DeskewCount
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_RANGE                  775:768
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_MSB                        775
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_LSB                        768
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_REL_RANGE              775:768
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_REL_MSB                    775
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_REL_LSB                    768
`define DCM_DESKEWTABLEDESC_FPS16DESKEWCOUNT_RESET_VALUE              8'h17

// macros with short names for field Dcm_DeskewTableDesc.fps16DeskewCount
`define DCM_DSKWTBLDSC_FPS16DSKWCNT_RANGE                           775:768
`define DCM_DSKWTBLDSC_FPS16DSKWCNT_MSB                                 775
`define DCM_DSKWTBLDSC_FPS16DSKWCNT_LSB                                 768
`define DCM_DSKWTBLDSC_FPS16DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS16DSKWCNT_RESET_VALUE                       8'h17

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps17DeskewCount
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_RANGE                  783:776
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_MSB                        783
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_LSB                        776
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_REL_RANGE              783:776
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_REL_MSB                    783
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_REL_LSB                    776
`define DCM_DESKEWTABLEDESC_FPS17DESKEWCOUNT_RESET_VALUE              8'h15

// macros with short names for field Dcm_DeskewTableDesc.fps17DeskewCount
`define DCM_DSKWTBLDSC_FPS17DSKWCNT_RANGE                           783:776
`define DCM_DSKWTBLDSC_FPS17DSKWCNT_MSB                                 783
`define DCM_DSKWTBLDSC_FPS17DSKWCNT_LSB                                 776
`define DCM_DSKWTBLDSC_FPS17DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS17DSKWCNT_RESET_VALUE                       8'h15

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps18DeskewCount
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_RANGE                  791:784
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_MSB                        791
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_LSB                        784
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_REL_RANGE              791:784
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_REL_MSB                    791
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_REL_LSB                    784
`define DCM_DESKEWTABLEDESC_FPS18DESKEWCOUNT_RESET_VALUE              8'h13

// macros with short names for field Dcm_DeskewTableDesc.fps18DeskewCount
`define DCM_DSKWTBLDSC_FPS18DSKWCNT_RANGE                           791:784
`define DCM_DSKWTBLDSC_FPS18DSKWCNT_MSB                                 791
`define DCM_DSKWTBLDSC_FPS18DSKWCNT_LSB                                 784
`define DCM_DSKWTBLDSC_FPS18DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS18DSKWCNT_RESET_VALUE                       8'h13

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps19DeskewCount
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_RANGE                  799:792
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_MSB                        799
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_LSB                        792
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_REL_RANGE              799:792
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_REL_MSB                    799
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_REL_LSB                    792
`define DCM_DESKEWTABLEDESC_FPS19DESKEWCOUNT_RESET_VALUE              8'h11

// macros with short names for field Dcm_DeskewTableDesc.fps19DeskewCount
`define DCM_DSKWTBLDSC_FPS19DSKWCNT_RANGE                           799:792
`define DCM_DSKWTBLDSC_FPS19DSKWCNT_MSB                                 799
`define DCM_DSKWTBLDSC_FPS19DSKWCNT_LSB                                 792
`define DCM_DSKWTBLDSC_FPS19DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS19DSKWCNT_RESET_VALUE                       8'h11

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps20DeskewCount
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_RANGE                  807:800
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_MSB                        807
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_LSB                        800
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_REL_RANGE              807:800
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_REL_MSB                    807
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_REL_LSB                    800
`define DCM_DESKEWTABLEDESC_FPS20DESKEWCOUNT_RESET_VALUE               8'hf

// macros with short names for field Dcm_DeskewTableDesc.fps20DeskewCount
`define DCM_DSKWTBLDSC_FPS20DSKWCNT_RANGE                           807:800
`define DCM_DSKWTBLDSC_FPS20DSKWCNT_MSB                                 807
`define DCM_DSKWTBLDSC_FPS20DSKWCNT_LSB                                 800
`define DCM_DSKWTBLDSC_FPS20DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS20DSKWCNT_RESET_VALUE                        8'hf

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps21DeskewCount
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_RANGE                  815:808
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_MSB                        815
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_LSB                        808
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_REL_RANGE              815:808
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_REL_MSB                    815
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_REL_LSB                    808
`define DCM_DESKEWTABLEDESC_FPS21DESKEWCOUNT_RESET_VALUE               8'hd

// macros with short names for field Dcm_DeskewTableDesc.fps21DeskewCount
`define DCM_DSKWTBLDSC_FPS21DSKWCNT_RANGE                           815:808
`define DCM_DSKWTBLDSC_FPS21DSKWCNT_MSB                                 815
`define DCM_DSKWTBLDSC_FPS21DSKWCNT_LSB                                 808
`define DCM_DSKWTBLDSC_FPS21DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS21DSKWCNT_RESET_VALUE                        8'hd

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps22DeskewCount
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_RANGE                  823:816
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_MSB                        823
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_LSB                        816
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_REL_RANGE              823:816
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_REL_MSB                    823
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_REL_LSB                    816
`define DCM_DESKEWTABLEDESC_FPS22DESKEWCOUNT_RESET_VALUE               8'hd

// macros with short names for field Dcm_DeskewTableDesc.fps22DeskewCount
`define DCM_DSKWTBLDSC_FPS22DSKWCNT_RANGE                           823:816
`define DCM_DSKWTBLDSC_FPS22DSKWCNT_MSB                                 823
`define DCM_DSKWTBLDSC_FPS22DSKWCNT_LSB                                 816
`define DCM_DSKWTBLDSC_FPS22DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS22DSKWCNT_RESET_VALUE                        8'hd

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps23DeskewCount
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_RANGE                  831:824
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_MSB                        831
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_LSB                        824
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_REL_RANGE              831:824
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_REL_MSB                    831
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_REL_LSB                    824
`define DCM_DESKEWTABLEDESC_FPS23DESKEWCOUNT_RESET_VALUE               8'hd

// macros with short names for field Dcm_DeskewTableDesc.fps23DeskewCount
`define DCM_DSKWTBLDSC_FPS23DSKWCNT_RANGE                           831:824
`define DCM_DSKWTBLDSC_FPS23DSKWCNT_MSB                                 831
`define DCM_DSKWTBLDSC_FPS23DSKWCNT_LSB                                 824
`define DCM_DSKWTBLDSC_FPS23DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS23DSKWCNT_RESET_VALUE                        8'hd

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.fps24DeskewCount
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_RANGE                  839:832
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_MSB                        839
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_LSB                        832
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_REL_RANGE              839:832
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_REL_MSB                    839
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_REL_LSB                    832
`define DCM_DESKEWTABLEDESC_FPS24DESKEWCOUNT_RESET_VALUE               8'hd

// macros with short names for field Dcm_DeskewTableDesc.fps24DeskewCount
`define DCM_DSKWTBLDSC_FPS24DSKWCNT_RANGE                           839:832
`define DCM_DSKWTBLDSC_FPS24DSKWCNT_MSB                                 839
`define DCM_DSKWTBLDSC_FPS24DSKWCNT_LSB                                 832
`define DCM_DSKWTBLDSC_FPS24DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_FPS24DSKWCNT_RESET_VALUE                        8'hd

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.egrDeskewCount
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_RANGE                    847:840
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_MSB                          847
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_LSB                          840
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_REL_RANGE                847:840
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_REL_MSB                      847
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_REL_LSB                      840
`define DCM_DESKEWTABLEDESC_EGRDESKEWCOUNT_RESET_VALUE                 8'hc

// macros with short names for field Dcm_DeskewTableDesc.egrDeskewCount
`define DCM_DSKWTBLDSC_EGRDSKWCNT_RANGE                             847:840
`define DCM_DSKWTBLDSC_EGRDSKWCNT_MSB                                   847
`define DCM_DSKWTBLDSC_EGRDSKWCNT_LSB                                   840
`define DCM_DSKWTBLDSC_EGRDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_EGRDSKWCNT_RESET_VALUE                          8'hc

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm17DeskewCount
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_RANGE                  855:848
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_MSB                        855
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_LSB                        848
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_WIDTH                        8
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_REL_RANGE              855:848
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_REL_MSB                    855
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_REL_LSB                    848
`define DCM_DESKEWTABLEDESC_DMM17DESKEWCOUNT_RESET_VALUE               8'h8

// macros with short names for field Dcm_DeskewTableDesc.dmm17DeskewCount
`define DCM_DSKWTBLDSC_DMM17DSKWCNT_RANGE                           855:848
`define DCM_DSKWTBLDSC_DMM17DSKWCNT_MSB                                 855
`define DCM_DSKWTBLDSC_DMM17DSKWCNT_LSB                                 848
`define DCM_DSKWTBLDSC_DMM17DSKWCNT_WIDTH                                 8
`define DCM_DSKWTBLDSC_DMM17DSKWCNT_RESET_VALUE                        8'h8

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.rweDeskewCount
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_RANGE                    863:856
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_MSB                          863
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_LSB                          856
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_REL_RANGE                863:856
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_REL_MSB                      863
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_REL_LSB                      856
`define DCM_DESKEWTABLEDESC_RWEDESKEWCOUNT_RESET_VALUE                 8'h9

// macros with short names for field Dcm_DeskewTableDesc.rweDeskewCount
`define DCM_DSKWTBLDSC_RWDSKWCNT_RANGE                              863:856
`define DCM_DSKWTBLDSC_RWDSKWCNT_MSB                                    863
`define DCM_DSKWTBLDSC_RWDSKWCNT_LSB                                    856
`define DCM_DSKWTBLDSC_RWDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_RWDSKWCNT_RESET_VALUE                           8'h9

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.epfDeskewCount
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_RANGE                    871:864
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_MSB                          871
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_LSB                          864
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_REL_RANGE                871:864
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_REL_MSB                      871
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_REL_LSB                      864
`define DCM_DESKEWTABLEDESC_EPFDESKEWCOUNT_RESET_VALUE                 8'h6

// macros with short names for field Dcm_DeskewTableDesc.epfDeskewCount
`define DCM_DSKWTBLDSC_EPFDSKWCNT_RANGE                             871:864
`define DCM_DSKWTBLDSC_EPFDSKWCNT_MSB                                   871
`define DCM_DSKWTBLDSC_EPFDSKWCNT_LSB                                   864
`define DCM_DSKWTBLDSC_EPFDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_EPFDSKWCNT_RESET_VALUE                          8'h6

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.dmm7DeskewCount
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_RANGE                   879:872
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_MSB                         879
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_LSB                         872
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_WIDTH                         8
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_REL_RANGE               879:872
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_REL_MSB                     879
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_REL_LSB                     872
`define DCM_DESKEWTABLEDESC_DMM7DESKEWCOUNT_RESET_VALUE                8'h3

// macros with short names for field Dcm_DeskewTableDesc.dmm7DeskewCount
`define DCM_DSKWTBLDSC_DMM7DSKWCNT_RANGE                            879:872
`define DCM_DSKWTBLDSC_DMM7DSKWCNT_MSB                                  879
`define DCM_DSKWTBLDSC_DMM7DSKWCNT_LSB                                  872
`define DCM_DSKWTBLDSC_DMM7DSKWCNT_WIDTH                                  8
`define DCM_DSKWTBLDSC_DMM7DSKWCNT_RESET_VALUE                         8'h3

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.mscEgressDeskewCount
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_RANGE              887:880
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_MSB                    887
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_LSB                    880
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_WIDTH                    8
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_REL_RANGE          887:880
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_REL_MSB                887
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_REL_LSB                880
`define DCM_DESKEWTABLEDESC_MSCEGRESSDESKEWCOUNT_RESET_VALUE           8'h2

// macros with short names for field Dcm_DeskewTableDesc.mscEgressDeskewCount
`define DCM_DSKWTBLDSC_MSCEGRSDSKWCNT_RANGE                         887:880
`define DCM_DSKWTBLDSC_MSCEGRSDSKWCNT_MSB                               887
`define DCM_DSKWTBLDSC_MSCEGRSDSKWCNT_LSB                               880
`define DCM_DSKWTBLDSC_MSCEGRSDSKWCNT_WIDTH                               8
`define DCM_DSKWTBLDSC_MSCEGRSDSKWCNT_RESET_VALUE                      8'h2

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.sliDeskewCount
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_RANGE                    895:888
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_MSB                          895
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_LSB                          888
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_REL_RANGE                895:888
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_REL_MSB                      895
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_REL_LSB                      888
`define DCM_DESKEWTABLEDESC_SLIDESKEWCOUNT_RESET_VALUE                8'hb4

// macros with short names for field Dcm_DeskewTableDesc.sliDeskewCount
`define DCM_DSKWTBLDSC_SLDSKWCNT_RANGE                              895:888
`define DCM_DSKWTBLDSC_SLDSKWCNT_MSB                                    895
`define DCM_DSKWTBLDSC_SLDSKWCNT_LSB                                    888
`define DCM_DSKWTBLDSC_SLDSKWCNT_WIDTH                                    8
`define DCM_DSKWTBLDSC_SLDSKWCNT_RESET_VALUE                          8'hb4

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_DeskewTableDesc.iqmDeskewCount
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_RANGE                    903:896
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_MSB                          903
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_LSB                          896
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_WIDTH                          8
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_REL_RANGE                903:896
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_REL_MSB                      903
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_REL_LSB                      896
`define DCM_DESKEWTABLEDESC_IQMDESKEWCOUNT_RESET_VALUE                8'h35

// macros with short names for field Dcm_DeskewTableDesc.iqmDeskewCount
`define DCM_DSKWTBLDSC_IQMDSKWCNT_RANGE                             903:896
`define DCM_DSKWTBLDSC_IQMDSKWCNT_MSB                                   903
`define DCM_DSKWTBLDSC_IQMDSKWCNT_LSB                                   896
`define DCM_DSKWTBLDSC_IQMDSKWCNT_WIDTH                                   8
`define DCM_DSKWTBLDSC_IQMDSKWCNT_RESET_VALUE                         8'h35

//macros for Register - Dcm_DeskewTableDesc
//Dcm_DeskewTableDesc is of type DcmDeskewTableDesc
`define DCM_DESKEWTABLEDESC_REG_NUM                                       1
`define DCM_DESKEWTABLEDESC_REG_ADDR                           32'h00000000
`define DCM_DESKEWTABLEDESC_REG_STRIDE                                  128
`define DCM_DESKEWTABLEDESC_REG_SIZE                                   1024
`define DCM_DESKEWTABLEDESC_REG_FPGA_NUM                                  0
`define DCM_DESKEWTABLEDESC_REG_PHY_SIZE                                904
`define DCM_DESKEWTABLEDESC_REG_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define DCM_DESKEWTABLEDESC_REG_ADDR_SIZE                                 0
`define DCM_DESKEWTABLEDESC_REG_RESET_VALUE xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx0011010110110100000000100000001100000110000010010000100000001100000011010000110100001101000011010000111100010001000100110001010100010111000110100001101100011110000111010010000100100000001000010010010100100100001001010010101000101001001011010010110100101111001100110011001100110101001101100011101000111011001111010011111101000001010000110100010101000111010010010100101101001101010011110101000101010011010101010101100001011001010110010101110101011100011000000110001001100001011000110110010001100110011010100110100101101100011011110110111101110000011100010111001001110011011101100111011101111000011110010111101001111100011111101000000010000000100000111000010110000111100010011000101110001101100011011000111110001111100100011001001110010101100101111001100110011011100111011001111110100001101000111010001110100011101001011010011110101001101010111010110110101110101100101011001110110100101101001011010110110110

// macros with short names for register Dcm_DeskewTableDesc
//Dcm_DeskewTableDesc is of type DcmDeskewTableDesc
`define DCM_DSKWTBLDSC_REG_NUM                                            1
`define DCM_DSKWTBLDSC_REG_ADDR                                32'h00000000
`define DCM_DSKWTBLDSC_REG_STRIDE                                       128
`define DCM_DSKWTBLDSC_REG_SIZE                                        1024
`define DCM_DSKWTBLDSC_REG_FPGA_NUM                                       0
`define DCM_DSKWTBLDSC_REG_PHY_SIZE                                     904

// macros for register Dcm_TlaIdTableDesc
//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.plcDcmId
`define DCM_TLAIDTABLEDESC_PLCDCMID_RANGE                               6:0
`define DCM_TLAIDTABLEDESC_PLCDCMID_MSB                                   6
`define DCM_TLAIDTABLEDESC_PLCDCMID_LSB                                   0
`define DCM_TLAIDTABLEDESC_PLCDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_PLCDCMID_REL_RANGE                           6:0
`define DCM_TLAIDTABLEDESC_PLCDCMID_REL_MSB                               6
`define DCM_TLAIDTABLEDESC_PLCDCMID_REL_LSB                               0
`define DCM_TLAIDTABLEDESC_PLCDCMID_RESET_VALUE                        7'h0

// macros with short names for field Dcm_TlaIdTableDesc.plcDcmId
`define DCM_TLIDTBLDSC_PLCDCMID_RANGE                                   6:0
`define DCM_TLIDTBLDSC_PLCDCMID_MSB                                       6
`define DCM_TLIDTBLDSC_PLCDCMID_LSB                                       0
`define DCM_TLIDTBLDSC_PLCDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_PLCDCMID_RESET_VALUE                            7'h0

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.nflDcmId
`define DCM_TLAIDTABLEDESC_NFLDCMID_RANGE                              13:7
`define DCM_TLAIDTABLEDESC_NFLDCMID_MSB                                  13
`define DCM_TLAIDTABLEDESC_NFLDCMID_LSB                                   7
`define DCM_TLAIDTABLEDESC_NFLDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NFLDCMID_REL_RANGE                          13:7
`define DCM_TLAIDTABLEDESC_NFLDCMID_REL_MSB                              13
`define DCM_TLAIDTABLEDESC_NFLDCMID_REL_LSB                               7
`define DCM_TLAIDTABLEDESC_NFLDCMID_RESET_VALUE                        7'h1

// macros with short names for field Dcm_TlaIdTableDesc.nflDcmId
`define DCM_TLIDTBLDSC_NFLDCMID_RANGE                                  13:7
`define DCM_TLIDTBLDSC_NFLDCMID_MSB                                      13
`define DCM_TLIDTBLDSC_NFLDCMID_LSB                                       7
`define DCM_TLIDTBLDSC_NFLDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_NFLDCMID_RESET_VALUE                            7'h1

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase0DcmId
`define DCM_TLAIDTABLEDESC_ASE0DCMID_RANGE                            20:14
`define DCM_TLAIDTABLEDESC_ASE0DCMID_MSB                                 20
`define DCM_TLAIDTABLEDESC_ASE0DCMID_LSB                                 14
`define DCM_TLAIDTABLEDESC_ASE0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE0DCMID_REL_RANGE                        20:14
`define DCM_TLAIDTABLEDESC_ASE0DCMID_REL_MSB                             20
`define DCM_TLAIDTABLEDESC_ASE0DCMID_REL_LSB                             14
`define DCM_TLAIDTABLEDESC_ASE0DCMID_RESET_VALUE                       7'h2

// macros with short names for field Dcm_TlaIdTableDesc.ase0DcmId
`define DCM_TLIDTBLDSC_AS0DCMID_RANGE                                 20:14
`define DCM_TLIDTBLDSC_AS0DCMID_MSB                                      20
`define DCM_TLIDTBLDSC_AS0DCMID_LSB                                      14
`define DCM_TLIDTBLDSC_AS0DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS0DCMID_RESET_VALUE                            7'h2

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase1DcmId
`define DCM_TLAIDTABLEDESC_ASE1DCMID_RANGE                            27:21
`define DCM_TLAIDTABLEDESC_ASE1DCMID_MSB                                 27
`define DCM_TLAIDTABLEDESC_ASE1DCMID_LSB                                 21
`define DCM_TLAIDTABLEDESC_ASE1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE1DCMID_REL_RANGE                        27:21
`define DCM_TLAIDTABLEDESC_ASE1DCMID_REL_MSB                             27
`define DCM_TLAIDTABLEDESC_ASE1DCMID_REL_LSB                             21
`define DCM_TLAIDTABLEDESC_ASE1DCMID_RESET_VALUE                       7'h3

// macros with short names for field Dcm_TlaIdTableDesc.ase1DcmId
`define DCM_TLIDTBLDSC_AS1DCMID_RANGE                                 27:21
`define DCM_TLIDTBLDSC_AS1DCMID_MSB                                      27
`define DCM_TLIDTBLDSC_AS1DCMID_LSB                                      21
`define DCM_TLIDTBLDSC_AS1DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS1DCMID_RESET_VALUE                            7'h3

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase2DcmId
`define DCM_TLAIDTABLEDESC_ASE2DCMID_RANGE                            34:28
`define DCM_TLAIDTABLEDESC_ASE2DCMID_MSB                                 34
`define DCM_TLAIDTABLEDESC_ASE2DCMID_LSB                                 28
`define DCM_TLAIDTABLEDESC_ASE2DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE2DCMID_REL_RANGE                        34:28
`define DCM_TLAIDTABLEDESC_ASE2DCMID_REL_MSB                             34
`define DCM_TLAIDTABLEDESC_ASE2DCMID_REL_LSB                             28
`define DCM_TLAIDTABLEDESC_ASE2DCMID_RESET_VALUE                       7'h4

// macros with short names for field Dcm_TlaIdTableDesc.ase2DcmId
`define DCM_TLIDTBLDSC_AS2DCMID_RANGE                                 34:28
`define DCM_TLIDTBLDSC_AS2DCMID_MSB                                      34
`define DCM_TLIDTBLDSC_AS2DCMID_LSB                                      28
`define DCM_TLIDTBLDSC_AS2DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS2DCMID_RESET_VALUE                            7'h4

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase3DcmId
`define DCM_TLAIDTABLEDESC_ASE3DCMID_RANGE                            41:35
`define DCM_TLAIDTABLEDESC_ASE3DCMID_MSB                                 41
`define DCM_TLAIDTABLEDESC_ASE3DCMID_LSB                                 35
`define DCM_TLAIDTABLEDESC_ASE3DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE3DCMID_REL_RANGE                        41:35
`define DCM_TLAIDTABLEDESC_ASE3DCMID_REL_MSB                             41
`define DCM_TLAIDTABLEDESC_ASE3DCMID_REL_LSB                             35
`define DCM_TLAIDTABLEDESC_ASE3DCMID_RESET_VALUE                       7'h5

// macros with short names for field Dcm_TlaIdTableDesc.ase3DcmId
`define DCM_TLIDTBLDSC_AS3DCMID_RANGE                                 41:35
`define DCM_TLIDTBLDSC_AS3DCMID_MSB                                      41
`define DCM_TLIDTBLDSC_AS3DCMID_LSB                                      35
`define DCM_TLIDTBLDSC_AS3DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS3DCMID_RESET_VALUE                            7'h5

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase4DcmId
`define DCM_TLAIDTABLEDESC_ASE4DCMID_RANGE                            48:42
`define DCM_TLAIDTABLEDESC_ASE4DCMID_MSB                                 48
`define DCM_TLAIDTABLEDESC_ASE4DCMID_LSB                                 42
`define DCM_TLAIDTABLEDESC_ASE4DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE4DCMID_REL_RANGE                        48:42
`define DCM_TLAIDTABLEDESC_ASE4DCMID_REL_MSB                             48
`define DCM_TLAIDTABLEDESC_ASE4DCMID_REL_LSB                             42
`define DCM_TLAIDTABLEDESC_ASE4DCMID_RESET_VALUE                       7'h6

// macros with short names for field Dcm_TlaIdTableDesc.ase4DcmId
`define DCM_TLIDTBLDSC_AS4DCMID_RANGE                                 48:42
`define DCM_TLIDTBLDSC_AS4DCMID_MSB                                      48
`define DCM_TLIDTBLDSC_AS4DCMID_LSB                                      42
`define DCM_TLIDTBLDSC_AS4DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS4DCMID_RESET_VALUE                            7'h6

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase5DcmId
`define DCM_TLAIDTABLEDESC_ASE5DCMID_RANGE                            55:49
`define DCM_TLAIDTABLEDESC_ASE5DCMID_MSB                                 55
`define DCM_TLAIDTABLEDESC_ASE5DCMID_LSB                                 49
`define DCM_TLAIDTABLEDESC_ASE5DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE5DCMID_REL_RANGE                        55:49
`define DCM_TLAIDTABLEDESC_ASE5DCMID_REL_MSB                             55
`define DCM_TLAIDTABLEDESC_ASE5DCMID_REL_LSB                             49
`define DCM_TLAIDTABLEDESC_ASE5DCMID_RESET_VALUE                       7'h7

// macros with short names for field Dcm_TlaIdTableDesc.ase5DcmId
`define DCM_TLIDTBLDSC_AS5DCMID_RANGE                                 55:49
`define DCM_TLIDTBLDSC_AS5DCMID_MSB                                      55
`define DCM_TLIDTBLDSC_AS5DCMID_LSB                                      49
`define DCM_TLIDTBLDSC_AS5DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS5DCMID_RESET_VALUE                            7'h7

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase6DcmId
`define DCM_TLAIDTABLEDESC_ASE6DCMID_RANGE                            62:56
`define DCM_TLAIDTABLEDESC_ASE6DCMID_MSB                                 62
`define DCM_TLAIDTABLEDESC_ASE6DCMID_LSB                                 56
`define DCM_TLAIDTABLEDESC_ASE6DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE6DCMID_REL_RANGE                        62:56
`define DCM_TLAIDTABLEDESC_ASE6DCMID_REL_MSB                             62
`define DCM_TLAIDTABLEDESC_ASE6DCMID_REL_LSB                             56
`define DCM_TLAIDTABLEDESC_ASE6DCMID_RESET_VALUE                       7'h8

// macros with short names for field Dcm_TlaIdTableDesc.ase6DcmId
`define DCM_TLIDTBLDSC_AS6DCMID_RANGE                                 62:56
`define DCM_TLIDTBLDSC_AS6DCMID_MSB                                      62
`define DCM_TLIDTBLDSC_AS6DCMID_LSB                                      56
`define DCM_TLIDTBLDSC_AS6DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS6DCMID_RESET_VALUE                            7'h8

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ase7DcmId
`define DCM_TLAIDTABLEDESC_ASE7DCMID_RANGE                            69:63
`define DCM_TLAIDTABLEDESC_ASE7DCMID_MSB                                 69
`define DCM_TLAIDTABLEDESC_ASE7DCMID_LSB                                 63
`define DCM_TLAIDTABLEDESC_ASE7DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_ASE7DCMID_REL_RANGE                        69:63
`define DCM_TLAIDTABLEDESC_ASE7DCMID_REL_MSB                             69
`define DCM_TLAIDTABLEDESC_ASE7DCMID_REL_LSB                             63
`define DCM_TLAIDTABLEDESC_ASE7DCMID_RESET_VALUE                       7'h9

// macros with short names for field Dcm_TlaIdTableDesc.ase7DcmId
`define DCM_TLIDTBLDSC_AS7DCMID_RANGE                                 69:63
`define DCM_TLIDTBLDSC_AS7DCMID_MSB                                      69
`define DCM_TLIDTBLDSC_AS7DCMID_LSB                                      63
`define DCM_TLIDTBLDSC_AS7DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AS7DCMID_RESET_VALUE                            7'h9

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.taq0DcmId
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_RANGE                            76:70
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_MSB                                 76
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_LSB                                 70
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_REL_RANGE                        76:70
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_REL_MSB                             76
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_REL_LSB                             70
`define DCM_TLAIDTABLEDESC_TAQ0DCMID_RESET_VALUE                       7'ha

// macros with short names for field Dcm_TlaIdTableDesc.taq0DcmId
`define DCM_TLIDTBLDSC_TQ0DCMID_RANGE                                 76:70
`define DCM_TLIDTBLDSC_TQ0DCMID_MSB                                      76
`define DCM_TLIDTBLDSC_TQ0DCMID_LSB                                      70
`define DCM_TLIDTBLDSC_TQ0DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TQ0DCMID_RESET_VALUE                            7'ha

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.taq1DcmId
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_RANGE                            83:77
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_MSB                                 83
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_LSB                                 77
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_REL_RANGE                        83:77
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_REL_MSB                             83
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_REL_LSB                             77
`define DCM_TLAIDTABLEDESC_TAQ1DCMID_RESET_VALUE                       7'hb

// macros with short names for field Dcm_TlaIdTableDesc.taq1DcmId
`define DCM_TLIDTBLDSC_TQ1DCMID_RANGE                                 83:77
`define DCM_TLIDTBLDSC_TQ1DCMID_MSB                                      83
`define DCM_TLIDTBLDSC_TQ1DCMID_LSB                                      77
`define DCM_TLIDTBLDSC_TQ1DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TQ1DCMID_RESET_VALUE                            7'hb

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.taq2DcmId
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_RANGE                            90:84
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_MSB                                 90
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_LSB                                 84
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_REL_RANGE                        90:84
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_REL_MSB                             90
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_REL_LSB                             84
`define DCM_TLAIDTABLEDESC_TAQ2DCMID_RESET_VALUE                       7'hc

// macros with short names for field Dcm_TlaIdTableDesc.taq2DcmId
`define DCM_TLIDTBLDSC_TQ2DCMID_RANGE                                 90:84
`define DCM_TLIDTBLDSC_TQ2DCMID_MSB                                      90
`define DCM_TLIDTBLDSC_TQ2DCMID_LSB                                      84
`define DCM_TLIDTBLDSC_TQ2DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TQ2DCMID_RESET_VALUE                            7'hc

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.taq3DcmId
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_RANGE                            97:91
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_MSB                                 97
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_LSB                                 91
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_REL_RANGE                        97:91
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_REL_MSB                             97
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_REL_LSB                             91
`define DCM_TLAIDTABLEDESC_TAQ3DCMID_RESET_VALUE                       7'hd

// macros with short names for field Dcm_TlaIdTableDesc.taq3DcmId
`define DCM_TLIDTBLDSC_TQ3DCMID_RANGE                                 97:91
`define DCM_TLIDTBLDSC_TQ3DCMID_MSB                                      97
`define DCM_TLIDTBLDSC_TQ3DCMID_LSB                                      91
`define DCM_TLIDTBLDSC_TQ3DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TQ3DCMID_RESET_VALUE                            7'hd

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.taq4DcmId
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_RANGE                           104:98
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_MSB                                104
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_LSB                                 98
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_REL_RANGE                       104:98
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_REL_MSB                            104
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_REL_LSB                             98
`define DCM_TLAIDTABLEDESC_TAQ4DCMID_RESET_VALUE                       7'he

// macros with short names for field Dcm_TlaIdTableDesc.taq4DcmId
`define DCM_TLIDTBLDSC_TQ4DCMID_RANGE                                104:98
`define DCM_TLIDTBLDSC_TQ4DCMID_MSB                                     104
`define DCM_TLIDTBLDSC_TQ4DCMID_LSB                                      98
`define DCM_TLIDTBLDSC_TQ4DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TQ4DCMID_RESET_VALUE                            7'he

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.taq5DcmId
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_RANGE                          111:105
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_MSB                                111
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_LSB                                105
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_REL_RANGE                      111:105
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_REL_MSB                            111
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_REL_LSB                            105
`define DCM_TLAIDTABLEDESC_TAQ5DCMID_RESET_VALUE                       7'hf

// macros with short names for field Dcm_TlaIdTableDesc.taq5DcmId
`define DCM_TLIDTBLDSC_TQ5DCMID_RANGE                               111:105
`define DCM_TLIDTBLDSC_TQ5DCMID_MSB                                     111
`define DCM_TLIDTBLDSC_TQ5DCMID_LSB                                     105
`define DCM_TLIDTBLDSC_TQ5DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TQ5DCMID_RESET_VALUE                            7'hf

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.taq6DcmId
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_RANGE                          118:112
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_MSB                                118
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_LSB                                112
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_REL_RANGE                      118:112
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_REL_MSB                            118
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_REL_LSB                            112
`define DCM_TLAIDTABLEDESC_TAQ6DCMID_RESET_VALUE                      7'h10

// macros with short names for field Dcm_TlaIdTableDesc.taq6DcmId
`define DCM_TLIDTBLDSC_TQ6DCMID_RANGE                               118:112
`define DCM_TLIDTBLDSC_TQ6DCMID_MSB                                     118
`define DCM_TLIDTBLDSC_TQ6DCMID_LSB                                     112
`define DCM_TLIDTBLDSC_TQ6DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TQ6DCMID_RESET_VALUE                           7'h10

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tlq0DcmId
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_RANGE                          125:119
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_MSB                                125
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_LSB                                119
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_REL_RANGE                      125:119
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_REL_MSB                            125
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_REL_LSB                            119
`define DCM_TLAIDTABLEDESC_TLQ0DCMID_RESET_VALUE                      7'h11

// macros with short names for field Dcm_TlaIdTableDesc.tlq0DcmId
`define DCM_TLIDTBLDSC_TLQ0DCMID_RANGE                              125:119
`define DCM_TLIDTBLDSC_TLQ0DCMID_MSB                                    125
`define DCM_TLIDTBLDSC_TLQ0DCMID_LSB                                    119
`define DCM_TLIDTBLDSC_TLQ0DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TLQ0DCMID_RESET_VALUE                          7'h11

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tlq1DcmId
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_RANGE                          132:126
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_MSB                                132
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_LSB                                126
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_REL_RANGE                      132:126
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_REL_MSB                            132
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_REL_LSB                            126
`define DCM_TLAIDTABLEDESC_TLQ1DCMID_RESET_VALUE                      7'h12

// macros with short names for field Dcm_TlaIdTableDesc.tlq1DcmId
`define DCM_TLIDTBLDSC_TLQ1DCMID_RANGE                              132:126
`define DCM_TLIDTBLDSC_TLQ1DCMID_MSB                                    132
`define DCM_TLIDTBLDSC_TLQ1DCMID_LSB                                    126
`define DCM_TLIDTBLDSC_TLQ1DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TLQ1DCMID_RESET_VALUE                          7'h12

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fse0DcmId
`define DCM_TLAIDTABLEDESC_FSE0DCMID_RANGE                          139:133
`define DCM_TLAIDTABLEDESC_FSE0DCMID_MSB                                139
`define DCM_TLAIDTABLEDESC_FSE0DCMID_LSB                                133
`define DCM_TLAIDTABLEDESC_FSE0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FSE0DCMID_REL_RANGE                      139:133
`define DCM_TLAIDTABLEDESC_FSE0DCMID_REL_MSB                            139
`define DCM_TLAIDTABLEDESC_FSE0DCMID_REL_LSB                            133
`define DCM_TLAIDTABLEDESC_FSE0DCMID_RESET_VALUE                      7'h13

// macros with short names for field Dcm_TlaIdTableDesc.fse0DcmId
`define DCM_TLIDTBLDSC_FS0DCMID_RANGE                               139:133
`define DCM_TLIDTBLDSC_FS0DCMID_MSB                                     139
`define DCM_TLIDTBLDSC_FS0DCMID_LSB                                     133
`define DCM_TLIDTBLDSC_FS0DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_FS0DCMID_RESET_VALUE                           7'h13

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fse1DcmId
`define DCM_TLAIDTABLEDESC_FSE1DCMID_RANGE                          146:140
`define DCM_TLAIDTABLEDESC_FSE1DCMID_MSB                                146
`define DCM_TLAIDTABLEDESC_FSE1DCMID_LSB                                140
`define DCM_TLAIDTABLEDESC_FSE1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FSE1DCMID_REL_RANGE                      146:140
`define DCM_TLAIDTABLEDESC_FSE1DCMID_REL_MSB                            146
`define DCM_TLAIDTABLEDESC_FSE1DCMID_REL_LSB                            140
`define DCM_TLAIDTABLEDESC_FSE1DCMID_RESET_VALUE                      7'h14

// macros with short names for field Dcm_TlaIdTableDesc.fse1DcmId
`define DCM_TLIDTBLDSC_FS1DCMID_RANGE                               146:140
`define DCM_TLIDTBLDSC_FS1DCMID_MSB                                     146
`define DCM_TLIDTBLDSC_FS1DCMID_LSB                                     140
`define DCM_TLIDTBLDSC_FS1DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_FS1DCMID_RESET_VALUE                           7'h14

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fse2DcmId
`define DCM_TLAIDTABLEDESC_FSE2DCMID_RANGE                          153:147
`define DCM_TLAIDTABLEDESC_FSE2DCMID_MSB                                153
`define DCM_TLAIDTABLEDESC_FSE2DCMID_LSB                                147
`define DCM_TLAIDTABLEDESC_FSE2DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FSE2DCMID_REL_RANGE                      153:147
`define DCM_TLAIDTABLEDESC_FSE2DCMID_REL_MSB                            153
`define DCM_TLAIDTABLEDESC_FSE2DCMID_REL_LSB                            147
`define DCM_TLAIDTABLEDESC_FSE2DCMID_RESET_VALUE                      7'h15

// macros with short names for field Dcm_TlaIdTableDesc.fse2DcmId
`define DCM_TLIDTBLDSC_FS2DCMID_RANGE                               153:147
`define DCM_TLIDTBLDSC_FS2DCMID_MSB                                     153
`define DCM_TLIDTBLDSC_FS2DCMID_LSB                                     147
`define DCM_TLIDTBLDSC_FS2DCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_FS2DCMID_RESET_VALUE                           7'h15

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.hsh0DcmId
`define DCM_TLAIDTABLEDESC_HSH0DCMID_RANGE                          160:154
`define DCM_TLAIDTABLEDESC_HSH0DCMID_MSB                                160
`define DCM_TLAIDTABLEDESC_HSH0DCMID_LSB                                154
`define DCM_TLAIDTABLEDESC_HSH0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_HSH0DCMID_REL_RANGE                      160:154
`define DCM_TLAIDTABLEDESC_HSH0DCMID_REL_MSB                            160
`define DCM_TLAIDTABLEDESC_HSH0DCMID_REL_LSB                            154
`define DCM_TLAIDTABLEDESC_HSH0DCMID_RESET_VALUE                      7'h16

// macros with short names for field Dcm_TlaIdTableDesc.hsh0DcmId
`define DCM_TLIDTBLDSC_HSH0DCMID_RANGE                              160:154
`define DCM_TLIDTBLDSC_HSH0DCMID_MSB                                    160
`define DCM_TLIDTBLDSC_HSH0DCMID_LSB                                    154
`define DCM_TLIDTBLDSC_HSH0DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_HSH0DCMID_RESET_VALUE                          7'h16

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.hsh1DcmId
`define DCM_TLAIDTABLEDESC_HSH1DCMID_RANGE                          167:161
`define DCM_TLAIDTABLEDESC_HSH1DCMID_MSB                                167
`define DCM_TLAIDTABLEDESC_HSH1DCMID_LSB                                161
`define DCM_TLAIDTABLEDESC_HSH1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_HSH1DCMID_REL_RANGE                      167:161
`define DCM_TLAIDTABLEDESC_HSH1DCMID_REL_MSB                            167
`define DCM_TLAIDTABLEDESC_HSH1DCMID_REL_LSB                            161
`define DCM_TLAIDTABLEDESC_HSH1DCMID_RESET_VALUE                      7'h17

// macros with short names for field Dcm_TlaIdTableDesc.hsh1DcmId
`define DCM_TLIDTBLDSC_HSH1DCMID_RANGE                              167:161
`define DCM_TLIDTBLDSC_HSH1DCMID_MSB                                    167
`define DCM_TLIDTBLDSC_HSH1DCMID_LSB                                    161
`define DCM_TLIDTBLDSC_HSH1DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_HSH1DCMID_RESET_VALUE                          7'h17

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.hsh2DcmId
`define DCM_TLAIDTABLEDESC_HSH2DCMID_RANGE                          174:168
`define DCM_TLAIDTABLEDESC_HSH2DCMID_MSB                                174
`define DCM_TLAIDTABLEDESC_HSH2DCMID_LSB                                168
`define DCM_TLAIDTABLEDESC_HSH2DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_HSH2DCMID_REL_RANGE                      174:168
`define DCM_TLAIDTABLEDESC_HSH2DCMID_REL_MSB                            174
`define DCM_TLAIDTABLEDESC_HSH2DCMID_REL_LSB                            168
`define DCM_TLAIDTABLEDESC_HSH2DCMID_RESET_VALUE                      7'h18

// macros with short names for field Dcm_TlaIdTableDesc.hsh2DcmId
`define DCM_TLIDTBLDSC_HSH2DCMID_RANGE                              174:168
`define DCM_TLIDTBLDSC_HSH2DCMID_MSB                                    174
`define DCM_TLIDTBLDSC_HSH2DCMID_LSB                                    168
`define DCM_TLIDTBLDSC_HSH2DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_HSH2DCMID_RESET_VALUE                          7'h18

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.hsh3DcmId
`define DCM_TLAIDTABLEDESC_HSH3DCMID_RANGE                          181:175
`define DCM_TLAIDTABLEDESC_HSH3DCMID_MSB                                181
`define DCM_TLAIDTABLEDESC_HSH3DCMID_LSB                                175
`define DCM_TLAIDTABLEDESC_HSH3DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_HSH3DCMID_REL_RANGE                      181:175
`define DCM_TLAIDTABLEDESC_HSH3DCMID_REL_MSB                            181
`define DCM_TLAIDTABLEDESC_HSH3DCMID_REL_LSB                            175
`define DCM_TLAIDTABLEDESC_HSH3DCMID_RESET_VALUE                      7'h19

// macros with short names for field Dcm_TlaIdTableDesc.hsh3DcmId
`define DCM_TLIDTBLDSC_HSH3DCMID_RANGE                              181:175
`define DCM_TLIDTBLDSC_HSH3DCMID_MSB                                    181
`define DCM_TLIDTBLDSC_HSH3DCMID_LSB                                    175
`define DCM_TLIDTBLDSC_HSH3DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_HSH3DCMID_RESET_VALUE                          7'h19

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.hsh4DcmId
`define DCM_TLAIDTABLEDESC_HSH4DCMID_RANGE                          188:182
`define DCM_TLAIDTABLEDESC_HSH4DCMID_MSB                                188
`define DCM_TLAIDTABLEDESC_HSH4DCMID_LSB                                182
`define DCM_TLAIDTABLEDESC_HSH4DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_HSH4DCMID_REL_RANGE                      188:182
`define DCM_TLAIDTABLEDESC_HSH4DCMID_REL_MSB                            188
`define DCM_TLAIDTABLEDESC_HSH4DCMID_REL_LSB                            182
`define DCM_TLAIDTABLEDESC_HSH4DCMID_RESET_VALUE                      7'h1a

// macros with short names for field Dcm_TlaIdTableDesc.hsh4DcmId
`define DCM_TLIDTBLDSC_HSH4DCMID_RANGE                              188:182
`define DCM_TLIDTBLDSC_HSH4DCMID_MSB                                    188
`define DCM_TLIDTBLDSC_HSH4DCMID_LSB                                    182
`define DCM_TLIDTBLDSC_HSH4DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_HSH4DCMID_RESET_VALUE                          7'h1a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.oft0DcmId
`define DCM_TLAIDTABLEDESC_OFT0DCMID_RANGE                          195:189
`define DCM_TLAIDTABLEDESC_OFT0DCMID_MSB                                195
`define DCM_TLAIDTABLEDESC_OFT0DCMID_LSB                                189
`define DCM_TLAIDTABLEDESC_OFT0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_OFT0DCMID_REL_RANGE                      195:189
`define DCM_TLAIDTABLEDESC_OFT0DCMID_REL_MSB                            195
`define DCM_TLAIDTABLEDESC_OFT0DCMID_REL_LSB                            189
`define DCM_TLAIDTABLEDESC_OFT0DCMID_RESET_VALUE                      7'h1b

// macros with short names for field Dcm_TlaIdTableDesc.oft0DcmId
`define DCM_TLIDTBLDSC_OFT0DCMID_RANGE                              195:189
`define DCM_TLIDTBLDSC_OFT0DCMID_MSB                                    195
`define DCM_TLIDTBLDSC_OFT0DCMID_LSB                                    189
`define DCM_TLIDTBLDSC_OFT0DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_OFT0DCMID_RESET_VALUE                          7'h1b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.oft1DcmId
`define DCM_TLAIDTABLEDESC_OFT1DCMID_RANGE                          202:196
`define DCM_TLAIDTABLEDESC_OFT1DCMID_MSB                                202
`define DCM_TLAIDTABLEDESC_OFT1DCMID_LSB                                196
`define DCM_TLAIDTABLEDESC_OFT1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_OFT1DCMID_REL_RANGE                      202:196
`define DCM_TLAIDTABLEDESC_OFT1DCMID_REL_MSB                            202
`define DCM_TLAIDTABLEDESC_OFT1DCMID_REL_LSB                            196
`define DCM_TLAIDTABLEDESC_OFT1DCMID_RESET_VALUE                      7'h1c

// macros with short names for field Dcm_TlaIdTableDesc.oft1DcmId
`define DCM_TLIDTBLDSC_OFT1DCMID_RANGE                              202:196
`define DCM_TLIDTBLDSC_OFT1DCMID_MSB                                    202
`define DCM_TLIDTBLDSC_OFT1DCMID_LSB                                    196
`define DCM_TLIDTBLDSC_OFT1DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_OFT1DCMID_RESET_VALUE                          7'h1c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tfq0DcmId
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_RANGE                          209:203
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_MSB                                209
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_LSB                                203
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_REL_RANGE                      209:203
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_REL_MSB                            209
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_REL_LSB                            203
`define DCM_TLAIDTABLEDESC_TFQ0DCMID_RESET_VALUE                      7'h1d

// macros with short names for field Dcm_TlaIdTableDesc.tfq0DcmId
`define DCM_TLIDTBLDSC_TFQ0DCMID_RANGE                              209:203
`define DCM_TLIDTBLDSC_TFQ0DCMID_MSB                                    209
`define DCM_TLIDTBLDSC_TFQ0DCMID_LSB                                    203
`define DCM_TLIDTBLDSC_TFQ0DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TFQ0DCMID_RESET_VALUE                          7'h1d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tfq1DcmId
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_RANGE                          216:210
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_MSB                                216
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_LSB                                210
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_REL_RANGE                      216:210
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_REL_MSB                            216
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_REL_LSB                            210
`define DCM_TLAIDTABLEDESC_TFQ1DCMID_RESET_VALUE                      7'h1e

// macros with short names for field Dcm_TlaIdTableDesc.tfq1DcmId
`define DCM_TLIDTBLDSC_TFQ1DCMID_RANGE                              216:210
`define DCM_TLIDTBLDSC_TFQ1DCMID_MSB                                    216
`define DCM_TLIDTBLDSC_TFQ1DCMID_LSB                                    210
`define DCM_TLIDTBLDSC_TFQ1DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TFQ1DCMID_RESET_VALUE                          7'h1e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.pimDcmId
`define DCM_TLAIDTABLEDESC_PIMDCMID_RANGE                           223:217
`define DCM_TLAIDTABLEDESC_PIMDCMID_MSB                                 223
`define DCM_TLAIDTABLEDESC_PIMDCMID_LSB                                 217
`define DCM_TLAIDTABLEDESC_PIMDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_PIMDCMID_REL_RANGE                       223:217
`define DCM_TLAIDTABLEDESC_PIMDCMID_REL_MSB                             223
`define DCM_TLAIDTABLEDESC_PIMDCMID_REL_LSB                             217
`define DCM_TLAIDTABLEDESC_PIMDCMID_RESET_VALUE                       7'h1f

// macros with short names for field Dcm_TlaIdTableDesc.pimDcmId
`define DCM_TLIDTBLDSC_PMDCMID_RANGE                                223:217
`define DCM_TLIDTBLDSC_PMDCMID_MSB                                      223
`define DCM_TLIDTBLDSC_PMDCMID_LSB                                      217
`define DCM_TLIDTBLDSC_PMDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_PMDCMID_RESET_VALUE                            7'h1f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.supDcmId
`define DCM_TLAIDTABLEDESC_SUPDCMID_RANGE                           230:224
`define DCM_TLAIDTABLEDESC_SUPDCMID_MSB                                 230
`define DCM_TLAIDTABLEDESC_SUPDCMID_LSB                                 224
`define DCM_TLAIDTABLEDESC_SUPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_SUPDCMID_REL_RANGE                       230:224
`define DCM_TLAIDTABLEDESC_SUPDCMID_REL_MSB                             230
`define DCM_TLAIDTABLEDESC_SUPDCMID_REL_LSB                             224
`define DCM_TLAIDTABLEDESC_SUPDCMID_RESET_VALUE                       7'h20

// macros with short names for field Dcm_TlaIdTableDesc.supDcmId
`define DCM_TLIDTBLDSC_SPDCMID_RANGE                                230:224
`define DCM_TLIDTBLDSC_SPDCMID_MSB                                      230
`define DCM_TLIDTBLDSC_SPDCMID_LSB                                      224
`define DCM_TLIDTBLDSC_SPDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_SPDCMID_RESET_VALUE                            7'h20

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.rmuDcmId
`define DCM_TLAIDTABLEDESC_RMUDCMID_RANGE                           237:231
`define DCM_TLAIDTABLEDESC_RMUDCMID_MSB                                 237
`define DCM_TLAIDTABLEDESC_RMUDCMID_LSB                                 231
`define DCM_TLAIDTABLEDESC_RMUDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_RMUDCMID_REL_RANGE                       237:231
`define DCM_TLAIDTABLEDESC_RMUDCMID_REL_MSB                             237
`define DCM_TLAIDTABLEDESC_RMUDCMID_REL_LSB                             231
`define DCM_TLAIDTABLEDESC_RMUDCMID_RESET_VALUE                       7'h21

// macros with short names for field Dcm_TlaIdTableDesc.rmuDcmId
`define DCM_TLIDTBLDSC_RMDCMID_RANGE                                237:231
`define DCM_TLIDTBLDSC_RMDCMID_MSB                                      237
`define DCM_TLIDTBLDSC_RMDCMID_LSB                                      231
`define DCM_TLIDTBLDSC_RMDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_RMDCMID_RESET_VALUE                            7'h21

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.secDcmId
`define DCM_TLAIDTABLEDESC_SECDCMID_RANGE                           244:238
`define DCM_TLAIDTABLEDESC_SECDCMID_MSB                                 244
`define DCM_TLAIDTABLEDESC_SECDCMID_LSB                                 238
`define DCM_TLAIDTABLEDESC_SECDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_SECDCMID_REL_RANGE                       244:238
`define DCM_TLAIDTABLEDESC_SECDCMID_REL_MSB                             244
`define DCM_TLAIDTABLEDESC_SECDCMID_REL_LSB                             238
`define DCM_TLAIDTABLEDESC_SECDCMID_RESET_VALUE                       7'h22

// macros with short names for field Dcm_TlaIdTableDesc.secDcmId
`define DCM_TLIDTBLDSC_SCDCMID_RANGE                                244:238
`define DCM_TLIDTBLDSC_SCDCMID_MSB                                      244
`define DCM_TLIDTBLDSC_SCDCMID_LSB                                      238
`define DCM_TLIDTBLDSC_SCDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_SCDCMID_RESET_VALUE                            7'h22

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.rreDcmId
`define DCM_TLAIDTABLEDESC_RREDCMID_RANGE                           251:245
`define DCM_TLAIDTABLEDESC_RREDCMID_MSB                                 251
`define DCM_TLAIDTABLEDESC_RREDCMID_LSB                                 245
`define DCM_TLAIDTABLEDESC_RREDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_RREDCMID_REL_RANGE                       251:245
`define DCM_TLAIDTABLEDESC_RREDCMID_REL_MSB                             251
`define DCM_TLAIDTABLEDESC_RREDCMID_REL_LSB                             245
`define DCM_TLAIDTABLEDESC_RREDCMID_RESET_VALUE                       7'h23

// macros with short names for field Dcm_TlaIdTableDesc.rreDcmId
`define DCM_TLIDTBLDSC_RRDCMID_RANGE                                251:245
`define DCM_TLIDTBLDSC_RRDCMID_MSB                                      251
`define DCM_TLIDTBLDSC_RRDCMID_LSB                                      245
`define DCM_TLIDTBLDSC_RRDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_RRDCMID_RESET_VALUE                            7'h23

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.nifDcmId
`define DCM_TLAIDTABLEDESC_NIFDCMID_RANGE                           258:252
`define DCM_TLAIDTABLEDESC_NIFDCMID_MSB                                 258
`define DCM_TLAIDTABLEDESC_NIFDCMID_LSB                                 252
`define DCM_TLAIDTABLEDESC_NIFDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NIFDCMID_REL_RANGE                       258:252
`define DCM_TLAIDTABLEDESC_NIFDCMID_REL_MSB                             258
`define DCM_TLAIDTABLEDESC_NIFDCMID_REL_LSB                             252
`define DCM_TLAIDTABLEDESC_NIFDCMID_RESET_VALUE                       7'h24

// macros with short names for field Dcm_TlaIdTableDesc.nifDcmId
`define DCM_TLIDTBLDSC_NFDCMID_RANGE                                258:252
`define DCM_TLIDTBLDSC_NFDCMID_MSB                                      258
`define DCM_TLIDTBLDSC_NFDCMID_LSB                                      252
`define DCM_TLIDTBLDSC_NFDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_NFDCMID_RESET_VALUE                            7'h24

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ipfDcmId
`define DCM_TLAIDTABLEDESC_IPFDCMID_RANGE                           265:259
`define DCM_TLAIDTABLEDESC_IPFDCMID_MSB                                 265
`define DCM_TLAIDTABLEDESC_IPFDCMID_LSB                                 259
`define DCM_TLAIDTABLEDESC_IPFDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_IPFDCMID_REL_RANGE                       265:259
`define DCM_TLAIDTABLEDESC_IPFDCMID_REL_MSB                             265
`define DCM_TLAIDTABLEDESC_IPFDCMID_REL_LSB                             259
`define DCM_TLAIDTABLEDESC_IPFDCMID_RESET_VALUE                       7'h25

// macros with short names for field Dcm_TlaIdTableDesc.ipfDcmId
`define DCM_TLIDTBLDSC_IPFDCMID_RANGE                               265:259
`define DCM_TLIDTBLDSC_IPFDCMID_MSB                                     265
`define DCM_TLIDTBLDSC_IPFDCMID_LSB                                     259
`define DCM_TLIDTBLDSC_IPFDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_IPFDCMID_RESET_VALUE                           7'h25

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fpeIngressDcmId
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_RANGE                    272:266
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_MSB                          272
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_LSB                          266
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_WIDTH                          7
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_REL_RANGE                272:266
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_REL_MSB                      272
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_REL_LSB                      266
`define DCM_TLAIDTABLEDESC_FPEINGRESSDCMID_RESET_VALUE                7'h26

// macros with short names for field Dcm_TlaIdTableDesc.fpeIngressDcmId
`define DCM_TLIDTBLDSC_FPINGRDCMID_RANGE                            272:266
`define DCM_TLIDTBLDSC_FPINGRDCMID_MSB                                  272
`define DCM_TLIDTBLDSC_FPINGRDCMID_LSB                                  266
`define DCM_TLIDTBLDSC_FPINGRDCMID_WIDTH                                  7
`define DCM_TLIDTBLDSC_FPINGRDCMID_RESET_VALUE                        7'h26

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fpeEgressDcmId
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_RANGE                     279:273
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_MSB                           279
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_LSB                           273
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_WIDTH                           7
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_REL_RANGE                 279:273
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_REL_MSB                       279
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_REL_LSB                       273
`define DCM_TLAIDTABLEDESC_FPEEGRESSDCMID_RESET_VALUE                 7'h27

// macros with short names for field Dcm_TlaIdTableDesc.fpeEgressDcmId
`define DCM_TLIDTBLDSC_FPEGRSDCMID_RANGE                            279:273
`define DCM_TLIDTBLDSC_FPEGRSDCMID_MSB                                  279
`define DCM_TLIDTBLDSC_FPEGRSDCMID_LSB                                  273
`define DCM_TLIDTBLDSC_FPEGRSDCMID_WIDTH                                  7
`define DCM_TLIDTBLDSC_FPEGRSDCMID_RESET_VALUE                        7'h27

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.cmmDcmId
`define DCM_TLAIDTABLEDESC_CMMDCMID_RANGE                           286:280
`define DCM_TLAIDTABLEDESC_CMMDCMID_MSB                                 286
`define DCM_TLAIDTABLEDESC_CMMDCMID_LSB                                 280
`define DCM_TLAIDTABLEDESC_CMMDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_CMMDCMID_REL_RANGE                       286:280
`define DCM_TLAIDTABLEDESC_CMMDCMID_REL_MSB                             286
`define DCM_TLAIDTABLEDESC_CMMDCMID_REL_LSB                             280
`define DCM_TLAIDTABLEDESC_CMMDCMID_RESET_VALUE                       7'h28

// macros with short names for field Dcm_TlaIdTableDesc.cmmDcmId
`define DCM_TLIDTBLDSC_CMMDCMID_RANGE                               286:280
`define DCM_TLIDTBLDSC_CMMDCMID_MSB                                     286
`define DCM_TLIDTBLDSC_CMMDCMID_LSB                                     280
`define DCM_TLIDTBLDSC_CMMDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_CMMDCMID_RESET_VALUE                           7'h28

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ippDcmId
`define DCM_TLAIDTABLEDESC_IPPDCMID_RANGE                           293:287
`define DCM_TLAIDTABLEDESC_IPPDCMID_MSB                                 293
`define DCM_TLAIDTABLEDESC_IPPDCMID_LSB                                 287
`define DCM_TLAIDTABLEDESC_IPPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_IPPDCMID_REL_RANGE                       293:287
`define DCM_TLAIDTABLEDESC_IPPDCMID_REL_MSB                             293
`define DCM_TLAIDTABLEDESC_IPPDCMID_REL_LSB                             287
`define DCM_TLAIDTABLEDESC_IPPDCMID_RESET_VALUE                       7'h29

// macros with short names for field Dcm_TlaIdTableDesc.ippDcmId
`define DCM_TLIDTBLDSC_IPPDCMID_RANGE                               293:287
`define DCM_TLIDTBLDSC_IPPDCMID_MSB                                     293
`define DCM_TLIDTBLDSC_IPPDCMID_LSB                                     287
`define DCM_TLIDTBLDSC_IPPDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_IPPDCMID_RESET_VALUE                           7'h29

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ileDcmId
`define DCM_TLAIDTABLEDESC_ILEDCMID_RANGE                           300:294
`define DCM_TLAIDTABLEDESC_ILEDCMID_MSB                                 300
`define DCM_TLAIDTABLEDESC_ILEDCMID_LSB                                 294
`define DCM_TLAIDTABLEDESC_ILEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_ILEDCMID_REL_RANGE                       300:294
`define DCM_TLAIDTABLEDESC_ILEDCMID_REL_MSB                             300
`define DCM_TLAIDTABLEDESC_ILEDCMID_REL_LSB                             294
`define DCM_TLAIDTABLEDESC_ILEDCMID_RESET_VALUE                       7'h2a

// macros with short names for field Dcm_TlaIdTableDesc.ileDcmId
`define DCM_TLIDTBLDSC_ILDCMID_RANGE                                300:294
`define DCM_TLIDTBLDSC_ILDCMID_MSB                                      300
`define DCM_TLIDTBLDSC_ILDCMID_LSB                                      294
`define DCM_TLIDTBLDSC_ILDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_ILDCMID_RESET_VALUE                            7'h2a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps0DcmId
`define DCM_TLAIDTABLEDESC_FPS0DCMID_RANGE                          307:301
`define DCM_TLAIDTABLEDESC_FPS0DCMID_MSB                                307
`define DCM_TLAIDTABLEDESC_FPS0DCMID_LSB                                301
`define DCM_TLAIDTABLEDESC_FPS0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS0DCMID_REL_RANGE                      307:301
`define DCM_TLAIDTABLEDESC_FPS0DCMID_REL_MSB                            307
`define DCM_TLAIDTABLEDESC_FPS0DCMID_REL_LSB                            301
`define DCM_TLAIDTABLEDESC_FPS0DCMID_RESET_VALUE                      7'h2b

// macros with short names for field Dcm_TlaIdTableDesc.fps0DcmId
`define DCM_TLIDTBLDSC_FPS0DCMID_RANGE                              307:301
`define DCM_TLIDTBLDSC_FPS0DCMID_MSB                                    307
`define DCM_TLIDTBLDSC_FPS0DCMID_LSB                                    301
`define DCM_TLIDTBLDSC_FPS0DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS0DCMID_RESET_VALUE                          7'h2b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps1DcmId
`define DCM_TLAIDTABLEDESC_FPS1DCMID_RANGE                          314:308
`define DCM_TLAIDTABLEDESC_FPS1DCMID_MSB                                314
`define DCM_TLAIDTABLEDESC_FPS1DCMID_LSB                                308
`define DCM_TLAIDTABLEDESC_FPS1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS1DCMID_REL_RANGE                      314:308
`define DCM_TLAIDTABLEDESC_FPS1DCMID_REL_MSB                            314
`define DCM_TLAIDTABLEDESC_FPS1DCMID_REL_LSB                            308
`define DCM_TLAIDTABLEDESC_FPS1DCMID_RESET_VALUE                      7'h2c

// macros with short names for field Dcm_TlaIdTableDesc.fps1DcmId
`define DCM_TLIDTBLDSC_FPS1DCMID_RANGE                              314:308
`define DCM_TLIDTBLDSC_FPS1DCMID_MSB                                    314
`define DCM_TLIDTBLDSC_FPS1DCMID_LSB                                    308
`define DCM_TLIDTBLDSC_FPS1DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS1DCMID_RESET_VALUE                          7'h2c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps2DcmId
`define DCM_TLAIDTABLEDESC_FPS2DCMID_RANGE                          321:315
`define DCM_TLAIDTABLEDESC_FPS2DCMID_MSB                                321
`define DCM_TLAIDTABLEDESC_FPS2DCMID_LSB                                315
`define DCM_TLAIDTABLEDESC_FPS2DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS2DCMID_REL_RANGE                      321:315
`define DCM_TLAIDTABLEDESC_FPS2DCMID_REL_MSB                            321
`define DCM_TLAIDTABLEDESC_FPS2DCMID_REL_LSB                            315
`define DCM_TLAIDTABLEDESC_FPS2DCMID_RESET_VALUE                      7'h2d

// macros with short names for field Dcm_TlaIdTableDesc.fps2DcmId
`define DCM_TLIDTBLDSC_FPS2DCMID_RANGE                              321:315
`define DCM_TLIDTBLDSC_FPS2DCMID_MSB                                    321
`define DCM_TLIDTBLDSC_FPS2DCMID_LSB                                    315
`define DCM_TLIDTBLDSC_FPS2DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS2DCMID_RESET_VALUE                          7'h2d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps3DcmId
`define DCM_TLAIDTABLEDESC_FPS3DCMID_RANGE                          328:322
`define DCM_TLAIDTABLEDESC_FPS3DCMID_MSB                                328
`define DCM_TLAIDTABLEDESC_FPS3DCMID_LSB                                322
`define DCM_TLAIDTABLEDESC_FPS3DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS3DCMID_REL_RANGE                      328:322
`define DCM_TLAIDTABLEDESC_FPS3DCMID_REL_MSB                            328
`define DCM_TLAIDTABLEDESC_FPS3DCMID_REL_LSB                            322
`define DCM_TLAIDTABLEDESC_FPS3DCMID_RESET_VALUE                      7'h2e

// macros with short names for field Dcm_TlaIdTableDesc.fps3DcmId
`define DCM_TLIDTBLDSC_FPS3DCMID_RANGE                              328:322
`define DCM_TLIDTBLDSC_FPS3DCMID_MSB                                    328
`define DCM_TLIDTBLDSC_FPS3DCMID_LSB                                    322
`define DCM_TLIDTBLDSC_FPS3DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS3DCMID_RESET_VALUE                          7'h2e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps4DcmId
`define DCM_TLAIDTABLEDESC_FPS4DCMID_RANGE                          335:329
`define DCM_TLAIDTABLEDESC_FPS4DCMID_MSB                                335
`define DCM_TLAIDTABLEDESC_FPS4DCMID_LSB                                329
`define DCM_TLAIDTABLEDESC_FPS4DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS4DCMID_REL_RANGE                      335:329
`define DCM_TLAIDTABLEDESC_FPS4DCMID_REL_MSB                            335
`define DCM_TLAIDTABLEDESC_FPS4DCMID_REL_LSB                            329
`define DCM_TLAIDTABLEDESC_FPS4DCMID_RESET_VALUE                      7'h2f

// macros with short names for field Dcm_TlaIdTableDesc.fps4DcmId
`define DCM_TLIDTBLDSC_FPS4DCMID_RANGE                              335:329
`define DCM_TLIDTBLDSC_FPS4DCMID_MSB                                    335
`define DCM_TLIDTBLDSC_FPS4DCMID_LSB                                    329
`define DCM_TLIDTBLDSC_FPS4DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS4DCMID_RESET_VALUE                          7'h2f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps5DcmId
`define DCM_TLAIDTABLEDESC_FPS5DCMID_RANGE                          342:336
`define DCM_TLAIDTABLEDESC_FPS5DCMID_MSB                                342
`define DCM_TLAIDTABLEDESC_FPS5DCMID_LSB                                336
`define DCM_TLAIDTABLEDESC_FPS5DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS5DCMID_REL_RANGE                      342:336
`define DCM_TLAIDTABLEDESC_FPS5DCMID_REL_MSB                            342
`define DCM_TLAIDTABLEDESC_FPS5DCMID_REL_LSB                            336
`define DCM_TLAIDTABLEDESC_FPS5DCMID_RESET_VALUE                      7'h30

// macros with short names for field Dcm_TlaIdTableDesc.fps5DcmId
`define DCM_TLIDTBLDSC_FPS5DCMID_RANGE                              342:336
`define DCM_TLIDTBLDSC_FPS5DCMID_MSB                                    342
`define DCM_TLIDTBLDSC_FPS5DCMID_LSB                                    336
`define DCM_TLIDTBLDSC_FPS5DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS5DCMID_RESET_VALUE                          7'h30

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps6DcmId
`define DCM_TLAIDTABLEDESC_FPS6DCMID_RANGE                          349:343
`define DCM_TLAIDTABLEDESC_FPS6DCMID_MSB                                349
`define DCM_TLAIDTABLEDESC_FPS6DCMID_LSB                                343
`define DCM_TLAIDTABLEDESC_FPS6DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS6DCMID_REL_RANGE                      349:343
`define DCM_TLAIDTABLEDESC_FPS6DCMID_REL_MSB                            349
`define DCM_TLAIDTABLEDESC_FPS6DCMID_REL_LSB                            343
`define DCM_TLAIDTABLEDESC_FPS6DCMID_RESET_VALUE                      7'h31

// macros with short names for field Dcm_TlaIdTableDesc.fps6DcmId
`define DCM_TLIDTBLDSC_FPS6DCMID_RANGE                              349:343
`define DCM_TLIDTBLDSC_FPS6DCMID_MSB                                    349
`define DCM_TLIDTBLDSC_FPS6DCMID_LSB                                    343
`define DCM_TLIDTBLDSC_FPS6DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS6DCMID_RESET_VALUE                          7'h31

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps7DcmId
`define DCM_TLAIDTABLEDESC_FPS7DCMID_RANGE                          356:350
`define DCM_TLAIDTABLEDESC_FPS7DCMID_MSB                                356
`define DCM_TLAIDTABLEDESC_FPS7DCMID_LSB                                350
`define DCM_TLAIDTABLEDESC_FPS7DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS7DCMID_REL_RANGE                      356:350
`define DCM_TLAIDTABLEDESC_FPS7DCMID_REL_MSB                            356
`define DCM_TLAIDTABLEDESC_FPS7DCMID_REL_LSB                            350
`define DCM_TLAIDTABLEDESC_FPS7DCMID_RESET_VALUE                      7'h32

// macros with short names for field Dcm_TlaIdTableDesc.fps7DcmId
`define DCM_TLIDTBLDSC_FPS7DCMID_RANGE                              356:350
`define DCM_TLIDTBLDSC_FPS7DCMID_MSB                                    356
`define DCM_TLIDTBLDSC_FPS7DCMID_LSB                                    350
`define DCM_TLIDTBLDSC_FPS7DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS7DCMID_RESET_VALUE                          7'h32

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps8DcmId
`define DCM_TLAIDTABLEDESC_FPS8DCMID_RANGE                          363:357
`define DCM_TLAIDTABLEDESC_FPS8DCMID_MSB                                363
`define DCM_TLAIDTABLEDESC_FPS8DCMID_LSB                                357
`define DCM_TLAIDTABLEDESC_FPS8DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS8DCMID_REL_RANGE                      363:357
`define DCM_TLAIDTABLEDESC_FPS8DCMID_REL_MSB                            363
`define DCM_TLAIDTABLEDESC_FPS8DCMID_REL_LSB                            357
`define DCM_TLAIDTABLEDESC_FPS8DCMID_RESET_VALUE                      7'h33

// macros with short names for field Dcm_TlaIdTableDesc.fps8DcmId
`define DCM_TLIDTBLDSC_FPS8DCMID_RANGE                              363:357
`define DCM_TLIDTBLDSC_FPS8DCMID_MSB                                    363
`define DCM_TLIDTBLDSC_FPS8DCMID_LSB                                    357
`define DCM_TLIDTBLDSC_FPS8DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS8DCMID_RESET_VALUE                          7'h33

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps9DcmId
`define DCM_TLAIDTABLEDESC_FPS9DCMID_RANGE                          370:364
`define DCM_TLAIDTABLEDESC_FPS9DCMID_MSB                                370
`define DCM_TLAIDTABLEDESC_FPS9DCMID_LSB                                364
`define DCM_TLAIDTABLEDESC_FPS9DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_FPS9DCMID_REL_RANGE                      370:364
`define DCM_TLAIDTABLEDESC_FPS9DCMID_REL_MSB                            370
`define DCM_TLAIDTABLEDESC_FPS9DCMID_REL_LSB                            364
`define DCM_TLAIDTABLEDESC_FPS9DCMID_RESET_VALUE                      7'h34

// macros with short names for field Dcm_TlaIdTableDesc.fps9DcmId
`define DCM_TLIDTBLDSC_FPS9DCMID_RANGE                              370:364
`define DCM_TLIDTBLDSC_FPS9DCMID_MSB                                    370
`define DCM_TLIDTBLDSC_FPS9DCMID_LSB                                    364
`define DCM_TLIDTBLDSC_FPS9DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_FPS9DCMID_RESET_VALUE                          7'h34

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps10DcmId
`define DCM_TLAIDTABLEDESC_FPS10DCMID_RANGE                         377:371
`define DCM_TLAIDTABLEDESC_FPS10DCMID_MSB                               377
`define DCM_TLAIDTABLEDESC_FPS10DCMID_LSB                               371
`define DCM_TLAIDTABLEDESC_FPS10DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS10DCMID_REL_RANGE                     377:371
`define DCM_TLAIDTABLEDESC_FPS10DCMID_REL_MSB                           377
`define DCM_TLAIDTABLEDESC_FPS10DCMID_REL_LSB                           371
`define DCM_TLAIDTABLEDESC_FPS10DCMID_RESET_VALUE                     7'h35

// macros with short names for field Dcm_TlaIdTableDesc.fps10DcmId
`define DCM_TLIDTBLDSC_FPS10DCMID_RANGE                             377:371
`define DCM_TLIDTBLDSC_FPS10DCMID_MSB                                   377
`define DCM_TLIDTBLDSC_FPS10DCMID_LSB                                   371
`define DCM_TLIDTBLDSC_FPS10DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS10DCMID_RESET_VALUE                         7'h35

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps11DcmId
`define DCM_TLAIDTABLEDESC_FPS11DCMID_RANGE                         384:378
`define DCM_TLAIDTABLEDESC_FPS11DCMID_MSB                               384
`define DCM_TLAIDTABLEDESC_FPS11DCMID_LSB                               378
`define DCM_TLAIDTABLEDESC_FPS11DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS11DCMID_REL_RANGE                     384:378
`define DCM_TLAIDTABLEDESC_FPS11DCMID_REL_MSB                           384
`define DCM_TLAIDTABLEDESC_FPS11DCMID_REL_LSB                           378
`define DCM_TLAIDTABLEDESC_FPS11DCMID_RESET_VALUE                     7'h36

// macros with short names for field Dcm_TlaIdTableDesc.fps11DcmId
`define DCM_TLIDTBLDSC_FPS11DCMID_RANGE                             384:378
`define DCM_TLIDTBLDSC_FPS11DCMID_MSB                                   384
`define DCM_TLIDTBLDSC_FPS11DCMID_LSB                                   378
`define DCM_TLIDTBLDSC_FPS11DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS11DCMID_RESET_VALUE                         7'h36

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps12DcmId
`define DCM_TLAIDTABLEDESC_FPS12DCMID_RANGE                         391:385
`define DCM_TLAIDTABLEDESC_FPS12DCMID_MSB                               391
`define DCM_TLAIDTABLEDESC_FPS12DCMID_LSB                               385
`define DCM_TLAIDTABLEDESC_FPS12DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS12DCMID_REL_RANGE                     391:385
`define DCM_TLAIDTABLEDESC_FPS12DCMID_REL_MSB                           391
`define DCM_TLAIDTABLEDESC_FPS12DCMID_REL_LSB                           385
`define DCM_TLAIDTABLEDESC_FPS12DCMID_RESET_VALUE                     7'h37

// macros with short names for field Dcm_TlaIdTableDesc.fps12DcmId
`define DCM_TLIDTBLDSC_FPS12DCMID_RANGE                             391:385
`define DCM_TLIDTBLDSC_FPS12DCMID_MSB                                   391
`define DCM_TLIDTBLDSC_FPS12DCMID_LSB                                   385
`define DCM_TLIDTBLDSC_FPS12DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS12DCMID_RESET_VALUE                         7'h37

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps13DcmId
`define DCM_TLAIDTABLEDESC_FPS13DCMID_RANGE                         398:392
`define DCM_TLAIDTABLEDESC_FPS13DCMID_MSB                               398
`define DCM_TLAIDTABLEDESC_FPS13DCMID_LSB                               392
`define DCM_TLAIDTABLEDESC_FPS13DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS13DCMID_REL_RANGE                     398:392
`define DCM_TLAIDTABLEDESC_FPS13DCMID_REL_MSB                           398
`define DCM_TLAIDTABLEDESC_FPS13DCMID_REL_LSB                           392
`define DCM_TLAIDTABLEDESC_FPS13DCMID_RESET_VALUE                     7'h38

// macros with short names for field Dcm_TlaIdTableDesc.fps13DcmId
`define DCM_TLIDTBLDSC_FPS13DCMID_RANGE                             398:392
`define DCM_TLIDTBLDSC_FPS13DCMID_MSB                                   398
`define DCM_TLIDTBLDSC_FPS13DCMID_LSB                                   392
`define DCM_TLIDTBLDSC_FPS13DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS13DCMID_RESET_VALUE                         7'h38

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps14DcmId
`define DCM_TLAIDTABLEDESC_FPS14DCMID_RANGE                         405:399
`define DCM_TLAIDTABLEDESC_FPS14DCMID_MSB                               405
`define DCM_TLAIDTABLEDESC_FPS14DCMID_LSB                               399
`define DCM_TLAIDTABLEDESC_FPS14DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS14DCMID_REL_RANGE                     405:399
`define DCM_TLAIDTABLEDESC_FPS14DCMID_REL_MSB                           405
`define DCM_TLAIDTABLEDESC_FPS14DCMID_REL_LSB                           399
`define DCM_TLAIDTABLEDESC_FPS14DCMID_RESET_VALUE                     7'h39

// macros with short names for field Dcm_TlaIdTableDesc.fps14DcmId
`define DCM_TLIDTBLDSC_FPS14DCMID_RANGE                             405:399
`define DCM_TLIDTBLDSC_FPS14DCMID_MSB                                   405
`define DCM_TLIDTBLDSC_FPS14DCMID_LSB                                   399
`define DCM_TLIDTBLDSC_FPS14DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS14DCMID_RESET_VALUE                         7'h39

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps15DcmId
`define DCM_TLAIDTABLEDESC_FPS15DCMID_RANGE                         412:406
`define DCM_TLAIDTABLEDESC_FPS15DCMID_MSB                               412
`define DCM_TLAIDTABLEDESC_FPS15DCMID_LSB                               406
`define DCM_TLAIDTABLEDESC_FPS15DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS15DCMID_REL_RANGE                     412:406
`define DCM_TLAIDTABLEDESC_FPS15DCMID_REL_MSB                           412
`define DCM_TLAIDTABLEDESC_FPS15DCMID_REL_LSB                           406
`define DCM_TLAIDTABLEDESC_FPS15DCMID_RESET_VALUE                     7'h3a

// macros with short names for field Dcm_TlaIdTableDesc.fps15DcmId
`define DCM_TLIDTBLDSC_FPS15DCMID_RANGE                             412:406
`define DCM_TLIDTBLDSC_FPS15DCMID_MSB                                   412
`define DCM_TLIDTBLDSC_FPS15DCMID_LSB                                   406
`define DCM_TLIDTBLDSC_FPS15DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS15DCMID_RESET_VALUE                         7'h3a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps16DcmId
`define DCM_TLAIDTABLEDESC_FPS16DCMID_RANGE                         419:413
`define DCM_TLAIDTABLEDESC_FPS16DCMID_MSB                               419
`define DCM_TLAIDTABLEDESC_FPS16DCMID_LSB                               413
`define DCM_TLAIDTABLEDESC_FPS16DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS16DCMID_REL_RANGE                     419:413
`define DCM_TLAIDTABLEDESC_FPS16DCMID_REL_MSB                           419
`define DCM_TLAIDTABLEDESC_FPS16DCMID_REL_LSB                           413
`define DCM_TLAIDTABLEDESC_FPS16DCMID_RESET_VALUE                     7'h3b

// macros with short names for field Dcm_TlaIdTableDesc.fps16DcmId
`define DCM_TLIDTBLDSC_FPS16DCMID_RANGE                             419:413
`define DCM_TLIDTBLDSC_FPS16DCMID_MSB                                   419
`define DCM_TLIDTBLDSC_FPS16DCMID_LSB                                   413
`define DCM_TLIDTBLDSC_FPS16DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS16DCMID_RESET_VALUE                         7'h3b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps17DcmId
`define DCM_TLAIDTABLEDESC_FPS17DCMID_RANGE                         426:420
`define DCM_TLAIDTABLEDESC_FPS17DCMID_MSB                               426
`define DCM_TLAIDTABLEDESC_FPS17DCMID_LSB                               420
`define DCM_TLAIDTABLEDESC_FPS17DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS17DCMID_REL_RANGE                     426:420
`define DCM_TLAIDTABLEDESC_FPS17DCMID_REL_MSB                           426
`define DCM_TLAIDTABLEDESC_FPS17DCMID_REL_LSB                           420
`define DCM_TLAIDTABLEDESC_FPS17DCMID_RESET_VALUE                     7'h3c

// macros with short names for field Dcm_TlaIdTableDesc.fps17DcmId
`define DCM_TLIDTBLDSC_FPS17DCMID_RANGE                             426:420
`define DCM_TLIDTBLDSC_FPS17DCMID_MSB                                   426
`define DCM_TLIDTBLDSC_FPS17DCMID_LSB                                   420
`define DCM_TLIDTBLDSC_FPS17DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS17DCMID_RESET_VALUE                         7'h3c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps18DcmId
`define DCM_TLAIDTABLEDESC_FPS18DCMID_RANGE                         433:427
`define DCM_TLAIDTABLEDESC_FPS18DCMID_MSB                               433
`define DCM_TLAIDTABLEDESC_FPS18DCMID_LSB                               427
`define DCM_TLAIDTABLEDESC_FPS18DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS18DCMID_REL_RANGE                     433:427
`define DCM_TLAIDTABLEDESC_FPS18DCMID_REL_MSB                           433
`define DCM_TLAIDTABLEDESC_FPS18DCMID_REL_LSB                           427
`define DCM_TLAIDTABLEDESC_FPS18DCMID_RESET_VALUE                     7'h3d

// macros with short names for field Dcm_TlaIdTableDesc.fps18DcmId
`define DCM_TLIDTBLDSC_FPS18DCMID_RANGE                             433:427
`define DCM_TLIDTBLDSC_FPS18DCMID_MSB                                   433
`define DCM_TLIDTBLDSC_FPS18DCMID_LSB                                   427
`define DCM_TLIDTBLDSC_FPS18DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS18DCMID_RESET_VALUE                         7'h3d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps19DcmId
`define DCM_TLAIDTABLEDESC_FPS19DCMID_RANGE                         440:434
`define DCM_TLAIDTABLEDESC_FPS19DCMID_MSB                               440
`define DCM_TLAIDTABLEDESC_FPS19DCMID_LSB                               434
`define DCM_TLAIDTABLEDESC_FPS19DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS19DCMID_REL_RANGE                     440:434
`define DCM_TLAIDTABLEDESC_FPS19DCMID_REL_MSB                           440
`define DCM_TLAIDTABLEDESC_FPS19DCMID_REL_LSB                           434
`define DCM_TLAIDTABLEDESC_FPS19DCMID_RESET_VALUE                     7'h3e

// macros with short names for field Dcm_TlaIdTableDesc.fps19DcmId
`define DCM_TLIDTBLDSC_FPS19DCMID_RANGE                             440:434
`define DCM_TLIDTBLDSC_FPS19DCMID_MSB                                   440
`define DCM_TLIDTBLDSC_FPS19DCMID_LSB                                   434
`define DCM_TLIDTBLDSC_FPS19DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS19DCMID_RESET_VALUE                         7'h3e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps20DcmId
`define DCM_TLAIDTABLEDESC_FPS20DCMID_RANGE                         447:441
`define DCM_TLAIDTABLEDESC_FPS20DCMID_MSB                               447
`define DCM_TLAIDTABLEDESC_FPS20DCMID_LSB                               441
`define DCM_TLAIDTABLEDESC_FPS20DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS20DCMID_REL_RANGE                     447:441
`define DCM_TLAIDTABLEDESC_FPS20DCMID_REL_MSB                           447
`define DCM_TLAIDTABLEDESC_FPS20DCMID_REL_LSB                           441
`define DCM_TLAIDTABLEDESC_FPS20DCMID_RESET_VALUE                     7'h3f

// macros with short names for field Dcm_TlaIdTableDesc.fps20DcmId
`define DCM_TLIDTBLDSC_FPS20DCMID_RANGE                             447:441
`define DCM_TLIDTBLDSC_FPS20DCMID_MSB                                   447
`define DCM_TLIDTBLDSC_FPS20DCMID_LSB                                   441
`define DCM_TLIDTBLDSC_FPS20DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS20DCMID_RESET_VALUE                         7'h3f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps21DcmId
`define DCM_TLAIDTABLEDESC_FPS21DCMID_RANGE                         454:448
`define DCM_TLAIDTABLEDESC_FPS21DCMID_MSB                               454
`define DCM_TLAIDTABLEDESC_FPS21DCMID_LSB                               448
`define DCM_TLAIDTABLEDESC_FPS21DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS21DCMID_REL_RANGE                     454:448
`define DCM_TLAIDTABLEDESC_FPS21DCMID_REL_MSB                           454
`define DCM_TLAIDTABLEDESC_FPS21DCMID_REL_LSB                           448
`define DCM_TLAIDTABLEDESC_FPS21DCMID_RESET_VALUE                     7'h40

// macros with short names for field Dcm_TlaIdTableDesc.fps21DcmId
`define DCM_TLIDTBLDSC_FPS21DCMID_RANGE                             454:448
`define DCM_TLIDTBLDSC_FPS21DCMID_MSB                                   454
`define DCM_TLIDTBLDSC_FPS21DCMID_LSB                                   448
`define DCM_TLIDTBLDSC_FPS21DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS21DCMID_RESET_VALUE                         7'h40

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps22DcmId
`define DCM_TLAIDTABLEDESC_FPS22DCMID_RANGE                         461:455
`define DCM_TLAIDTABLEDESC_FPS22DCMID_MSB                               461
`define DCM_TLAIDTABLEDESC_FPS22DCMID_LSB                               455
`define DCM_TLAIDTABLEDESC_FPS22DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS22DCMID_REL_RANGE                     461:455
`define DCM_TLAIDTABLEDESC_FPS22DCMID_REL_MSB                           461
`define DCM_TLAIDTABLEDESC_FPS22DCMID_REL_LSB                           455
`define DCM_TLAIDTABLEDESC_FPS22DCMID_RESET_VALUE                     7'h41

// macros with short names for field Dcm_TlaIdTableDesc.fps22DcmId
`define DCM_TLIDTBLDSC_FPS22DCMID_RANGE                             461:455
`define DCM_TLIDTBLDSC_FPS22DCMID_MSB                                   461
`define DCM_TLIDTBLDSC_FPS22DCMID_LSB                                   455
`define DCM_TLIDTBLDSC_FPS22DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS22DCMID_RESET_VALUE                         7'h41

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps23DcmId
`define DCM_TLAIDTABLEDESC_FPS23DCMID_RANGE                         468:462
`define DCM_TLAIDTABLEDESC_FPS23DCMID_MSB                               468
`define DCM_TLAIDTABLEDESC_FPS23DCMID_LSB                               462
`define DCM_TLAIDTABLEDESC_FPS23DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS23DCMID_REL_RANGE                     468:462
`define DCM_TLAIDTABLEDESC_FPS23DCMID_REL_MSB                           468
`define DCM_TLAIDTABLEDESC_FPS23DCMID_REL_LSB                           462
`define DCM_TLAIDTABLEDESC_FPS23DCMID_RESET_VALUE                     7'h42

// macros with short names for field Dcm_TlaIdTableDesc.fps23DcmId
`define DCM_TLIDTBLDSC_FPS23DCMID_RANGE                             468:462
`define DCM_TLIDTBLDSC_FPS23DCMID_MSB                                   468
`define DCM_TLIDTBLDSC_FPS23DCMID_LSB                                   462
`define DCM_TLIDTBLDSC_FPS23DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS23DCMID_RESET_VALUE                         7'h42

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fps24DcmId
`define DCM_TLAIDTABLEDESC_FPS24DCMID_RANGE                         475:469
`define DCM_TLAIDTABLEDESC_FPS24DCMID_MSB                               475
`define DCM_TLAIDTABLEDESC_FPS24DCMID_LSB                               469
`define DCM_TLAIDTABLEDESC_FPS24DCMID_WIDTH                               7
`define DCM_TLAIDTABLEDESC_FPS24DCMID_REL_RANGE                     475:469
`define DCM_TLAIDTABLEDESC_FPS24DCMID_REL_MSB                           475
`define DCM_TLAIDTABLEDESC_FPS24DCMID_REL_LSB                           469
`define DCM_TLAIDTABLEDESC_FPS24DCMID_RESET_VALUE                     7'h43

// macros with short names for field Dcm_TlaIdTableDesc.fps24DcmId
`define DCM_TLIDTBLDSC_FPS24DCMID_RANGE                             475:469
`define DCM_TLIDTBLDSC_FPS24DCMID_MSB                                   475
`define DCM_TLIDTBLDSC_FPS24DCMID_LSB                                   469
`define DCM_TLIDTBLDSC_FPS24DCMID_WIDTH                                   7
`define DCM_TLIDTBLDSC_FPS24DCMID_RESET_VALUE                         7'h43

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.igrDcmId
`define DCM_TLAIDTABLEDESC_IGRDCMID_RANGE                           482:476
`define DCM_TLAIDTABLEDESC_IGRDCMID_MSB                                 482
`define DCM_TLAIDTABLEDESC_IGRDCMID_LSB                                 476
`define DCM_TLAIDTABLEDESC_IGRDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_IGRDCMID_REL_RANGE                       482:476
`define DCM_TLAIDTABLEDESC_IGRDCMID_REL_MSB                             482
`define DCM_TLAIDTABLEDESC_IGRDCMID_REL_LSB                             476
`define DCM_TLAIDTABLEDESC_IGRDCMID_RESET_VALUE                       7'h44

// macros with short names for field Dcm_TlaIdTableDesc.igrDcmId
`define DCM_TLIDTBLDSC_IGRDCMID_RANGE                               482:476
`define DCM_TLIDTBLDSC_IGRDCMID_MSB                                     482
`define DCM_TLIDTBLDSC_IGRDCMID_LSB                                     476
`define DCM_TLIDTBLDSC_IGRDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_IGRDCMID_RESET_VALUE                           7'h44

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.iqsDcmId
`define DCM_TLAIDTABLEDESC_IQSDCMID_RANGE                           489:483
`define DCM_TLAIDTABLEDESC_IQSDCMID_MSB                                 489
`define DCM_TLAIDTABLEDESC_IQSDCMID_LSB                                 483
`define DCM_TLAIDTABLEDESC_IQSDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_IQSDCMID_REL_RANGE                       489:483
`define DCM_TLAIDTABLEDESC_IQSDCMID_REL_MSB                             489
`define DCM_TLAIDTABLEDESC_IQSDCMID_REL_LSB                             483
`define DCM_TLAIDTABLEDESC_IQSDCMID_RESET_VALUE                       7'h45

// macros with short names for field Dcm_TlaIdTableDesc.iqsDcmId
`define DCM_TLIDTBLDSC_IQSDCMID_RANGE                               489:483
`define DCM_TLIDTBLDSC_IQSDCMID_MSB                                     489
`define DCM_TLIDTBLDSC_IQSDCMID_LSB                                     483
`define DCM_TLIDTBLDSC_IQSDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_IQSDCMID_RESET_VALUE                           7'h45

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.sqsDcmId
`define DCM_TLAIDTABLEDESC_SQSDCMID_RANGE                           496:490
`define DCM_TLAIDTABLEDESC_SQSDCMID_MSB                                 496
`define DCM_TLAIDTABLEDESC_SQSDCMID_LSB                                 490
`define DCM_TLAIDTABLEDESC_SQSDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_SQSDCMID_REL_RANGE                       496:490
`define DCM_TLAIDTABLEDESC_SQSDCMID_REL_MSB                             496
`define DCM_TLAIDTABLEDESC_SQSDCMID_REL_LSB                             490
`define DCM_TLAIDTABLEDESC_SQSDCMID_RESET_VALUE                       7'h46

// macros with short names for field Dcm_TlaIdTableDesc.sqsDcmId
`define DCM_TLIDTBLDSC_SQSDCMID_RANGE                               496:490
`define DCM_TLIDTBLDSC_SQSDCMID_MSB                                     496
`define DCM_TLIDTBLDSC_SQSDCMID_LSB                                     490
`define DCM_TLIDTBLDSC_SQSDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_SQSDCMID_RESET_VALUE                           7'h46

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.aqmDcmId
`define DCM_TLAIDTABLEDESC_AQMDCMID_RANGE                           503:497
`define DCM_TLAIDTABLEDESC_AQMDCMID_MSB                                 503
`define DCM_TLAIDTABLEDESC_AQMDCMID_LSB                                 497
`define DCM_TLAIDTABLEDESC_AQMDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_AQMDCMID_REL_RANGE                       503:497
`define DCM_TLAIDTABLEDESC_AQMDCMID_REL_MSB                             503
`define DCM_TLAIDTABLEDESC_AQMDCMID_REL_LSB                             497
`define DCM_TLAIDTABLEDESC_AQMDCMID_RESET_VALUE                       7'h47

// macros with short names for field Dcm_TlaIdTableDesc.aqmDcmId
`define DCM_TLIDTBLDSC_AQMDCMID_RANGE                               503:497
`define DCM_TLIDTBLDSC_AQMDCMID_MSB                                     503
`define DCM_TLIDTBLDSC_AQMDCMID_LSB                                     497
`define DCM_TLIDTBLDSC_AQMDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_AQMDCMID_RESET_VALUE                           7'h47

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.eqcDcmId
`define DCM_TLAIDTABLEDESC_EQCDCMID_RANGE                           510:504
`define DCM_TLAIDTABLEDESC_EQCDCMID_MSB                                 510
`define DCM_TLAIDTABLEDESC_EQCDCMID_LSB                                 504
`define DCM_TLAIDTABLEDESC_EQCDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_EQCDCMID_REL_RANGE                       510:504
`define DCM_TLAIDTABLEDESC_EQCDCMID_REL_MSB                             510
`define DCM_TLAIDTABLEDESC_EQCDCMID_REL_LSB                             504
`define DCM_TLAIDTABLEDESC_EQCDCMID_RESET_VALUE                       7'h48

// macros with short names for field Dcm_TlaIdTableDesc.eqcDcmId
`define DCM_TLIDTBLDSC_EQCDCMID_RANGE                               510:504
`define DCM_TLIDTBLDSC_EQCDCMID_MSB                                     510
`define DCM_TLIDTBLDSC_EQCDCMID_LSB                                     504
`define DCM_TLIDTBLDSC_EQCDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_EQCDCMID_RESET_VALUE                           7'h48

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.esmDcmId
`define DCM_TLAIDTABLEDESC_ESMDCMID_RANGE                           517:511
`define DCM_TLAIDTABLEDESC_ESMDCMID_MSB                                 517
`define DCM_TLAIDTABLEDESC_ESMDCMID_LSB                                 511
`define DCM_TLAIDTABLEDESC_ESMDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_ESMDCMID_REL_RANGE                       517:511
`define DCM_TLAIDTABLEDESC_ESMDCMID_REL_MSB                             517
`define DCM_TLAIDTABLEDESC_ESMDCMID_REL_LSB                             511
`define DCM_TLAIDTABLEDESC_ESMDCMID_RESET_VALUE                       7'h49

// macros with short names for field Dcm_TlaIdTableDesc.esmDcmId
`define DCM_TLIDTBLDSC_ESMDCMID_RANGE                               517:511
`define DCM_TLIDTBLDSC_ESMDCMID_MSB                                     517
`define DCM_TLIDTBLDSC_ESMDCMID_LSB                                     511
`define DCM_TLIDTBLDSC_ESMDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_ESMDCMID_RESET_VALUE                           7'h49

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.pbcDcmId
`define DCM_TLAIDTABLEDESC_PBCDCMID_RANGE                           524:518
`define DCM_TLAIDTABLEDESC_PBCDCMID_MSB                                 524
`define DCM_TLAIDTABLEDESC_PBCDCMID_LSB                                 518
`define DCM_TLAIDTABLEDESC_PBCDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_PBCDCMID_REL_RANGE                       524:518
`define DCM_TLAIDTABLEDESC_PBCDCMID_REL_MSB                             524
`define DCM_TLAIDTABLEDESC_PBCDCMID_REL_LSB                             518
`define DCM_TLAIDTABLEDESC_PBCDCMID_RESET_VALUE                       7'h4a

// macros with short names for field Dcm_TlaIdTableDesc.pbcDcmId
`define DCM_TLIDTBLDSC_PBCDCMID_RANGE                               524:518
`define DCM_TLIDTBLDSC_PBCDCMID_MSB                                     524
`define DCM_TLIDTBLDSC_PBCDCMID_LSB                                     518
`define DCM_TLIDTBLDSC_PBCDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_PBCDCMID_RESET_VALUE                           7'h4a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.sifDcmId
`define DCM_TLAIDTABLEDESC_SIFDCMID_RANGE                           531:525
`define DCM_TLAIDTABLEDESC_SIFDCMID_MSB                                 531
`define DCM_TLAIDTABLEDESC_SIFDCMID_LSB                                 525
`define DCM_TLAIDTABLEDESC_SIFDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_SIFDCMID_REL_RANGE                       531:525
`define DCM_TLAIDTABLEDESC_SIFDCMID_REL_MSB                             531
`define DCM_TLAIDTABLEDESC_SIFDCMID_REL_LSB                             525
`define DCM_TLAIDTABLEDESC_SIFDCMID_RESET_VALUE                       7'h4b

// macros with short names for field Dcm_TlaIdTableDesc.sifDcmId
`define DCM_TLIDTBLDSC_SFDCMID_RANGE                                531:525
`define DCM_TLIDTBLDSC_SFDCMID_MSB                                      531
`define DCM_TLIDTBLDSC_SFDCMID_LSB                                      525
`define DCM_TLIDTBLDSC_SFDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_SFDCMID_RESET_VALUE                            7'h4b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.frwDcmId
`define DCM_TLAIDTABLEDESC_FRWDCMID_RANGE                           538:532
`define DCM_TLAIDTABLEDESC_FRWDCMID_MSB                                 538
`define DCM_TLAIDTABLEDESC_FRWDCMID_LSB                                 532
`define DCM_TLAIDTABLEDESC_FRWDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_FRWDCMID_REL_RANGE                       538:532
`define DCM_TLAIDTABLEDESC_FRWDCMID_REL_MSB                             538
`define DCM_TLAIDTABLEDESC_FRWDCMID_REL_LSB                             532
`define DCM_TLAIDTABLEDESC_FRWDCMID_RESET_VALUE                       7'h4c

// macros with short names for field Dcm_TlaIdTableDesc.frwDcmId
`define DCM_TLIDTBLDSC_FRWDCMID_RANGE                               538:532
`define DCM_TLIDTBLDSC_FRWDCMID_MSB                                     538
`define DCM_TLIDTBLDSC_FRWDCMID_LSB                                     532
`define DCM_TLIDTBLDSC_FRWDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_FRWDCMID_RESET_VALUE                           7'h4c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.eppDcmId
`define DCM_TLAIDTABLEDESC_EPPDCMID_RANGE                           545:539
`define DCM_TLAIDTABLEDESC_EPPDCMID_MSB                                 545
`define DCM_TLAIDTABLEDESC_EPPDCMID_LSB                                 539
`define DCM_TLAIDTABLEDESC_EPPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_EPPDCMID_REL_RANGE                       545:539
`define DCM_TLAIDTABLEDESC_EPPDCMID_REL_MSB                             545
`define DCM_TLAIDTABLEDESC_EPPDCMID_REL_LSB                             539
`define DCM_TLAIDTABLEDESC_EPPDCMID_RESET_VALUE                       7'h4d

// macros with short names for field Dcm_TlaIdTableDesc.eppDcmId
`define DCM_TLIDTBLDSC_EPPDCMID_RANGE                               545:539
`define DCM_TLIDTBLDSC_EPPDCMID_MSB                                     545
`define DCM_TLIDTBLDSC_EPPDCMID_LSB                                     539
`define DCM_TLIDTBLDSC_EPPDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_EPPDCMID_RESET_VALUE                           7'h4d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.eleDcmId
`define DCM_TLAIDTABLEDESC_ELEDCMID_RANGE                           552:546
`define DCM_TLAIDTABLEDESC_ELEDCMID_MSB                                 552
`define DCM_TLAIDTABLEDESC_ELEDCMID_LSB                                 546
`define DCM_TLAIDTABLEDESC_ELEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_ELEDCMID_REL_RANGE                       552:546
`define DCM_TLAIDTABLEDESC_ELEDCMID_REL_MSB                             552
`define DCM_TLAIDTABLEDESC_ELEDCMID_REL_LSB                             546
`define DCM_TLAIDTABLEDESC_ELEDCMID_RESET_VALUE                       7'h4e

// macros with short names for field Dcm_TlaIdTableDesc.eleDcmId
`define DCM_TLIDTBLDSC_ELDCMID_RANGE                                552:546
`define DCM_TLIDTBLDSC_ELDCMID_MSB                                      552
`define DCM_TLIDTBLDSC_ELDCMID_LSB                                      546
`define DCM_TLIDTBLDSC_ELDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_ELDCMID_RESET_VALUE                            7'h4e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.egrDcmId
`define DCM_TLAIDTABLEDESC_EGRDCMID_RANGE                           559:553
`define DCM_TLAIDTABLEDESC_EGRDCMID_MSB                                 559
`define DCM_TLAIDTABLEDESC_EGRDCMID_LSB                                 553
`define DCM_TLAIDTABLEDESC_EGRDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_EGRDCMID_REL_RANGE                       559:553
`define DCM_TLAIDTABLEDESC_EGRDCMID_REL_MSB                             559
`define DCM_TLAIDTABLEDESC_EGRDCMID_REL_LSB                             553
`define DCM_TLAIDTABLEDESC_EGRDCMID_RESET_VALUE                       7'h4f

// macros with short names for field Dcm_TlaIdTableDesc.egrDcmId
`define DCM_TLIDTBLDSC_EGRDCMID_RANGE                               559:553
`define DCM_TLIDTBLDSC_EGRDCMID_MSB                                     559
`define DCM_TLIDTBLDSC_EGRDCMID_LSB                                     553
`define DCM_TLIDTBLDSC_EGRDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_EGRDCMID_RESET_VALUE                           7'h4f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.rweDcmId
`define DCM_TLAIDTABLEDESC_RWEDCMID_RANGE                           566:560
`define DCM_TLAIDTABLEDESC_RWEDCMID_MSB                                 566
`define DCM_TLAIDTABLEDESC_RWEDCMID_LSB                                 560
`define DCM_TLAIDTABLEDESC_RWEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_RWEDCMID_REL_RANGE                       566:560
`define DCM_TLAIDTABLEDESC_RWEDCMID_REL_MSB                             566
`define DCM_TLAIDTABLEDESC_RWEDCMID_REL_LSB                             560
`define DCM_TLAIDTABLEDESC_RWEDCMID_RESET_VALUE                       7'h50

// macros with short names for field Dcm_TlaIdTableDesc.rweDcmId
`define DCM_TLIDTBLDSC_RWDCMID_RANGE                                566:560
`define DCM_TLIDTBLDSC_RWDCMID_MSB                                      566
`define DCM_TLIDTBLDSC_RWDCMID_LSB                                      560
`define DCM_TLIDTBLDSC_RWDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_RWDCMID_RESET_VALUE                            7'h50

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.epfDcmId
`define DCM_TLAIDTABLEDESC_EPFDCMID_RANGE                           573:567
`define DCM_TLAIDTABLEDESC_EPFDCMID_MSB                                 573
`define DCM_TLAIDTABLEDESC_EPFDCMID_LSB                                 567
`define DCM_TLAIDTABLEDESC_EPFDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_EPFDCMID_REL_RANGE                       573:567
`define DCM_TLAIDTABLEDESC_EPFDCMID_REL_MSB                             573
`define DCM_TLAIDTABLEDESC_EPFDCMID_REL_LSB                             567
`define DCM_TLAIDTABLEDESC_EPFDCMID_RESET_VALUE                       7'h51

// macros with short names for field Dcm_TlaIdTableDesc.epfDcmId
`define DCM_TLIDTBLDSC_EPFDCMID_RANGE                               573:567
`define DCM_TLIDTBLDSC_EPFDCMID_MSB                                     573
`define DCM_TLIDTBLDSC_EPFDCMID_LSB                                     567
`define DCM_TLIDTBLDSC_EPFDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_EPFDCMID_RESET_VALUE                           7'h51

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.mscIngressDcmId
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_RANGE                    580:574
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_MSB                          580
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_LSB                          574
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_WIDTH                          7
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_REL_RANGE                580:574
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_REL_MSB                      580
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_REL_LSB                      574
`define DCM_TLAIDTABLEDESC_MSCINGRESSDCMID_RESET_VALUE                7'h52

// macros with short names for field Dcm_TlaIdTableDesc.mscIngressDcmId
`define DCM_TLIDTBLDSC_MSCINGRDCMID_RANGE                           580:574
`define DCM_TLIDTBLDSC_MSCINGRDCMID_MSB                                 580
`define DCM_TLIDTBLDSC_MSCINGRDCMID_LSB                                 574
`define DCM_TLIDTBLDSC_MSCINGRDCMID_WIDTH                                 7
`define DCM_TLIDTBLDSC_MSCINGRDCMID_RESET_VALUE                       7'h52

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.mscEgressDcmId
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_RANGE                     587:581
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_MSB                           587
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_LSB                           581
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_WIDTH                           7
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_REL_RANGE                 587:581
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_REL_MSB                       587
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_REL_LSB                       581
`define DCM_TLAIDTABLEDESC_MSCEGRESSDCMID_RESET_VALUE                 7'h53

// macros with short names for field Dcm_TlaIdTableDesc.mscEgressDcmId
`define DCM_TLIDTBLDSC_MSCEGRSDCMID_RANGE                           587:581
`define DCM_TLIDTBLDSC_MSCEGRSDCMID_MSB                                 587
`define DCM_TLIDTBLDSC_MSCEGRSDCMID_LSB                                 581
`define DCM_TLIDTBLDSC_MSCEGRSDCMID_WIDTH                                 7
`define DCM_TLIDTBLDSC_MSCEGRSDCMID_RESET_VALUE                       7'h53

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tsq0DcmId
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_RANGE                          594:588
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_MSB                                594
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_LSB                                588
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_REL_RANGE                      594:588
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_REL_MSB                            594
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_REL_LSB                            588
`define DCM_TLAIDTABLEDESC_TSQ0DCMID_RESET_VALUE                      7'h54

// macros with short names for field Dcm_TlaIdTableDesc.tsq0DcmId
`define DCM_TLIDTBLDSC_TSQ0DCMID_RANGE                              594:588
`define DCM_TLIDTBLDSC_TSQ0DCMID_MSB                                    594
`define DCM_TLIDTBLDSC_TSQ0DCMID_LSB                                    588
`define DCM_TLIDTBLDSC_TSQ0DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TSQ0DCMID_RESET_VALUE                          7'h54

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tsq1DcmId
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_RANGE                          601:595
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_MSB                                601
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_LSB                                595
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_REL_RANGE                      601:595
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_REL_MSB                            601
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_REL_LSB                            595
`define DCM_TLAIDTABLEDESC_TSQ1DCMID_RESET_VALUE                      7'h55

// macros with short names for field Dcm_TlaIdTableDesc.tsq1DcmId
`define DCM_TLIDTBLDSC_TSQ1DCMID_RANGE                              601:595
`define DCM_TLIDTBLDSC_TSQ1DCMID_MSB                                    601
`define DCM_TLIDTBLDSC_TSQ1DCMID_LSB                                    595
`define DCM_TLIDTBLDSC_TSQ1DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TSQ1DCMID_RESET_VALUE                          7'h55

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tsq2DcmId
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_RANGE                          608:602
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_MSB                                608
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_LSB                                602
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_REL_RANGE                      608:602
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_REL_MSB                            608
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_REL_LSB                            602
`define DCM_TLAIDTABLEDESC_TSQ2DCMID_RESET_VALUE                      7'h56

// macros with short names for field Dcm_TlaIdTableDesc.tsq2DcmId
`define DCM_TLIDTBLDSC_TSQ2DCMID_RANGE                              608:602
`define DCM_TLIDTBLDSC_TSQ2DCMID_MSB                                    608
`define DCM_TLIDTBLDSC_TSQ2DCMID_LSB                                    602
`define DCM_TLIDTBLDSC_TSQ2DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TSQ2DCMID_RESET_VALUE                          7'h56

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tsq3DcmId
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_RANGE                          615:609
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_MSB                                615
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_LSB                                609
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_WIDTH                                7
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_REL_RANGE                      615:609
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_REL_MSB                            615
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_REL_LSB                            609
`define DCM_TLAIDTABLEDESC_TSQ3DCMID_RESET_VALUE                      7'h57

// macros with short names for field Dcm_TlaIdTableDesc.tsq3DcmId
`define DCM_TLIDTBLDSC_TSQ3DCMID_RANGE                              615:609
`define DCM_TLIDTBLDSC_TSQ3DCMID_MSB                                    615
`define DCM_TLIDTBLDSC_TSQ3DCMID_LSB                                    609
`define DCM_TLIDTBLDSC_TSQ3DCMID_WIDTH                                    7
`define DCM_TLIDTBLDSC_TSQ3DCMID_RESET_VALUE                          7'h57

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.sliDcmId
`define DCM_TLAIDTABLEDESC_SLIDCMID_RANGE                           622:616
`define DCM_TLAIDTABLEDESC_SLIDCMID_MSB                                 622
`define DCM_TLAIDTABLEDESC_SLIDCMID_LSB                                 616
`define DCM_TLAIDTABLEDESC_SLIDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_SLIDCMID_REL_RANGE                       622:616
`define DCM_TLAIDTABLEDESC_SLIDCMID_REL_MSB                             622
`define DCM_TLAIDTABLEDESC_SLIDCMID_REL_LSB                             616
`define DCM_TLAIDTABLEDESC_SLIDCMID_RESET_VALUE                       7'h58

// macros with short names for field Dcm_TlaIdTableDesc.sliDcmId
`define DCM_TLIDTBLDSC_SLDCMID_RANGE                                622:616
`define DCM_TLIDTBLDSC_SLDCMID_MSB                                      622
`define DCM_TLIDTBLDSC_SLDCMID_LSB                                      616
`define DCM_TLIDTBLDSC_SLDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_SLDCMID_RESET_VALUE                            7'h58

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.iqmDcmId
`define DCM_TLAIDTABLEDESC_IQMDCMID_RANGE                           629:623
`define DCM_TLAIDTABLEDESC_IQMDCMID_MSB                                 629
`define DCM_TLAIDTABLEDESC_IQMDCMID_LSB                                 623
`define DCM_TLAIDTABLEDESC_IQMDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_IQMDCMID_REL_RANGE                       629:623
`define DCM_TLAIDTABLEDESC_IQMDCMID_REL_MSB                             629
`define DCM_TLAIDTABLEDESC_IQMDCMID_REL_LSB                             623
`define DCM_TLAIDTABLEDESC_IQMDCMID_RESET_VALUE                       7'h59

// macros with short names for field Dcm_TlaIdTableDesc.iqmDcmId
`define DCM_TLIDTBLDSC_IQMDCMID_RANGE                               629:623
`define DCM_TLIDTBLDSC_IQMDCMID_MSB                                     629
`define DCM_TLIDTBLDSC_IQMDCMID_LSB                                     623
`define DCM_TLIDTBLDSC_IQMDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_IQMDCMID_RESET_VALUE                           7'h59

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ismDcmId
`define DCM_TLAIDTABLEDESC_ISMDCMID_RANGE                           636:630
`define DCM_TLAIDTABLEDESC_ISMDCMID_MSB                                 636
`define DCM_TLAIDTABLEDESC_ISMDCMID_LSB                                 630
`define DCM_TLAIDTABLEDESC_ISMDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_ISMDCMID_REL_RANGE                       636:630
`define DCM_TLAIDTABLEDESC_ISMDCMID_REL_MSB                             636
`define DCM_TLAIDTABLEDESC_ISMDCMID_REL_LSB                             630
`define DCM_TLAIDTABLEDESC_ISMDCMID_RESET_VALUE                       7'h5a

// macros with short names for field Dcm_TlaIdTableDesc.ismDcmId
`define DCM_TLIDTBLDSC_ISMDCMID_RANGE                               636:630
`define DCM_TLIDTBLDSC_ISMDCMID_MSB                                     636
`define DCM_TLIDTBLDSC_ISMDCMID_LSB                                     630
`define DCM_TLIDTBLDSC_ISMDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_ISMDCMID_RESET_VALUE                           7'h5a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ftnDcmId
`define DCM_TLAIDTABLEDESC_FTNDCMID_RANGE                           643:637
`define DCM_TLAIDTABLEDESC_FTNDCMID_MSB                                 643
`define DCM_TLAIDTABLEDESC_FTNDCMID_LSB                                 637
`define DCM_TLAIDTABLEDESC_FTNDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_FTNDCMID_REL_RANGE                       643:637
`define DCM_TLAIDTABLEDESC_FTNDCMID_REL_MSB                             643
`define DCM_TLAIDTABLEDESC_FTNDCMID_REL_LSB                             637
`define DCM_TLAIDTABLEDESC_FTNDCMID_RESET_VALUE                       7'h5b

// macros with short names for field Dcm_TlaIdTableDesc.ftnDcmId
`define DCM_TLIDTBLDSC_FTNDCMID_RANGE                               643:637
`define DCM_TLIDTBLDSC_FTNDCMID_MSB                                     643
`define DCM_TLIDTBLDSC_FTNDCMID_LSB                                     637
`define DCM_TLIDTBLDSC_FTNDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_FTNDCMID_RESET_VALUE                           7'h5b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.svnDcmId
`define DCM_TLAIDTABLEDESC_SVNDCMID_RANGE                           650:644
`define DCM_TLAIDTABLEDESC_SVNDCMID_MSB                                 650
`define DCM_TLAIDTABLEDESC_SVNDCMID_LSB                                 644
`define DCM_TLAIDTABLEDESC_SVNDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_SVNDCMID_REL_RANGE                       650:644
`define DCM_TLAIDTABLEDESC_SVNDCMID_REL_MSB                             650
`define DCM_TLAIDTABLEDESC_SVNDCMID_REL_LSB                             644
`define DCM_TLAIDTABLEDESC_SVNDCMID_RESET_VALUE                       7'h5c

// macros with short names for field Dcm_TlaIdTableDesc.svnDcmId
`define DCM_TLIDTBLDSC_SVNDCMID_RANGE                               650:644
`define DCM_TLIDTBLDSC_SVNDCMID_MSB                                     650
`define DCM_TLIDTBLDSC_SVNDCMID_LSB                                     644
`define DCM_TLIDTBLDSC_SVNDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_SVNDCMID_RESET_VALUE                           7'h5c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.cciDcmId
`define DCM_TLAIDTABLEDESC_CCIDCMID_RANGE                           657:651
`define DCM_TLAIDTABLEDESC_CCIDCMID_MSB                                 657
`define DCM_TLAIDTABLEDESC_CCIDCMID_LSB                                 651
`define DCM_TLAIDTABLEDESC_CCIDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_CCIDCMID_REL_RANGE                       657:651
`define DCM_TLAIDTABLEDESC_CCIDCMID_REL_MSB                             657
`define DCM_TLAIDTABLEDESC_CCIDCMID_REL_LSB                             651
`define DCM_TLAIDTABLEDESC_CCIDCMID_RESET_VALUE                       7'h5d

// macros with short names for field Dcm_TlaIdTableDesc.cciDcmId
`define DCM_TLIDTBLDSC_CCDCMID_RANGE                                657:651
`define DCM_TLIDTBLDSC_CCDCMID_MSB                                      657
`define DCM_TLIDTBLDSC_CCDCMID_LSB                                      651
`define DCM_TLIDTBLDSC_CCDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_CCDCMID_RESET_VALUE                            7'h5d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.idtDcmId
`define DCM_TLAIDTABLEDESC_IDTDCMID_RANGE                           664:658
`define DCM_TLAIDTABLEDESC_IDTDCMID_MSB                                 664
`define DCM_TLAIDTABLEDESC_IDTDCMID_LSB                                 658
`define DCM_TLAIDTABLEDESC_IDTDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_IDTDCMID_REL_RANGE                       664:658
`define DCM_TLAIDTABLEDESC_IDTDCMID_REL_MSB                             664
`define DCM_TLAIDTABLEDESC_IDTDCMID_REL_LSB                             658
`define DCM_TLAIDTABLEDESC_IDTDCMID_RESET_VALUE                       7'h5e

// macros with short names for field Dcm_TlaIdTableDesc.idtDcmId
`define DCM_TLIDTBLDSC_IDTDCMID_RANGE                               664:658
`define DCM_TLIDTBLDSC_IDTDCMID_MSB                                     664
`define DCM_TLIDTBLDSC_IDTDCMID_LSB                                     658
`define DCM_TLIDTBLDSC_IDTDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_IDTDCMID_RESET_VALUE                           7'h5e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.napDcmId
`define DCM_TLAIDTABLEDESC_NAPDCMID_RANGE                           671:665
`define DCM_TLAIDTABLEDESC_NAPDCMID_MSB                                 671
`define DCM_TLAIDTABLEDESC_NAPDCMID_LSB                                 665
`define DCM_TLAIDTABLEDESC_NAPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NAPDCMID_REL_RANGE                       671:665
`define DCM_TLAIDTABLEDESC_NAPDCMID_REL_MSB                             671
`define DCM_TLAIDTABLEDESC_NAPDCMID_REL_LSB                             665
`define DCM_TLAIDTABLEDESC_NAPDCMID_RESET_VALUE                       7'h5f

// macros with short names for field Dcm_TlaIdTableDesc.napDcmId
`define DCM_TLIDTBLDSC_NPDCMID_RANGE                                671:665
`define DCM_TLIDTBLDSC_NPDCMID_MSB                                      671
`define DCM_TLIDTBLDSC_NPDCMID_LSB                                      665
`define DCM_TLIDTBLDSC_NPDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_NPDCMID_RESET_VALUE                            7'h5f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.treDcmId
`define DCM_TLAIDTABLEDESC_TREDCMID_RANGE                           678:672
`define DCM_TLAIDTABLEDESC_TREDCMID_MSB                                 678
`define DCM_TLAIDTABLEDESC_TREDCMID_LSB                                 672
`define DCM_TLAIDTABLEDESC_TREDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_TREDCMID_REL_RANGE                       678:672
`define DCM_TLAIDTABLEDESC_TREDCMID_REL_MSB                             678
`define DCM_TLAIDTABLEDESC_TREDCMID_REL_LSB                             672
`define DCM_TLAIDTABLEDESC_TREDCMID_RESET_VALUE                       7'h60

// macros with short names for field Dcm_TlaIdTableDesc.treDcmId
`define DCM_TLIDTBLDSC_TRDCMID_RANGE                                678:672
`define DCM_TLIDTBLDSC_TRDCMID_MSB                                      678
`define DCM_TLIDTBLDSC_TRDCMID_LSB                                      672
`define DCM_TLIDTBLDSC_TRDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_TRDCMID_RESET_VALUE                            7'h60

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ncbDcmId
`define DCM_TLAIDTABLEDESC_NCBDCMID_RANGE                           685:679
`define DCM_TLAIDTABLEDESC_NCBDCMID_MSB                                 685
`define DCM_TLAIDTABLEDESC_NCBDCMID_LSB                                 679
`define DCM_TLAIDTABLEDESC_NCBDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NCBDCMID_REL_RANGE                       685:679
`define DCM_TLAIDTABLEDESC_NCBDCMID_REL_MSB                             685
`define DCM_TLAIDTABLEDESC_NCBDCMID_REL_LSB                             679
`define DCM_TLAIDTABLEDESC_NCBDCMID_RESET_VALUE                       7'h61

// macros with short names for field Dcm_TlaIdTableDesc.ncbDcmId
`define DCM_TLIDTBLDSC_NCBDCMID_RANGE                               685:679
`define DCM_TLIDTBLDSC_NCBDCMID_MSB                                     685
`define DCM_TLIDTBLDSC_NCBDCMID_LSB                                     679
`define DCM_TLIDTBLDSC_NCBDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_NCBDCMID_RESET_VALUE                           7'h61

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.dpeDcmId
`define DCM_TLAIDTABLEDESC_DPEDCMID_RANGE                           692:686
`define DCM_TLAIDTABLEDESC_DPEDCMID_MSB                                 692
`define DCM_TLAIDTABLEDESC_DPEDCMID_LSB                                 686
`define DCM_TLAIDTABLEDESC_DPEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_DPEDCMID_REL_RANGE                       692:686
`define DCM_TLAIDTABLEDESC_DPEDCMID_REL_MSB                             692
`define DCM_TLAIDTABLEDESC_DPEDCMID_REL_LSB                             686
`define DCM_TLAIDTABLEDESC_DPEDCMID_RESET_VALUE                       7'h62

// macros with short names for field Dcm_TlaIdTableDesc.dpeDcmId
`define DCM_TLIDTBLDSC_DPDCMID_RANGE                                692:686
`define DCM_TLIDTBLDSC_DPDCMID_MSB                                      692
`define DCM_TLIDTBLDSC_DPDCMID_LSB                                      686
`define DCM_TLIDTBLDSC_DPDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_DPDCMID_RESET_VALUE                            7'h62

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.mceDcmId
`define DCM_TLAIDTABLEDESC_MCEDCMID_RANGE                           699:693
`define DCM_TLAIDTABLEDESC_MCEDCMID_MSB                                 699
`define DCM_TLAIDTABLEDESC_MCEDCMID_LSB                                 693
`define DCM_TLAIDTABLEDESC_MCEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_MCEDCMID_REL_RANGE                       699:693
`define DCM_TLAIDTABLEDESC_MCEDCMID_REL_MSB                             699
`define DCM_TLAIDTABLEDESC_MCEDCMID_REL_LSB                             693
`define DCM_TLAIDTABLEDESC_MCEDCMID_RESET_VALUE                       7'h63

// macros with short names for field Dcm_TlaIdTableDesc.mceDcmId
`define DCM_TLIDTBLDSC_MCDCMID_RANGE                                699:693
`define DCM_TLIDTBLDSC_MCDCMID_MSB                                      699
`define DCM_TLIDTBLDSC_MCDCMID_LSB                                      693
`define DCM_TLIDTBLDSC_MCDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_MCDCMID_RESET_VALUE                            7'h63

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.lkeDcmId
`define DCM_TLAIDTABLEDESC_LKEDCMID_RANGE                           706:700
`define DCM_TLAIDTABLEDESC_LKEDCMID_MSB                                 706
`define DCM_TLAIDTABLEDESC_LKEDCMID_LSB                                 700
`define DCM_TLAIDTABLEDESC_LKEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_LKEDCMID_REL_RANGE                       706:700
`define DCM_TLAIDTABLEDESC_LKEDCMID_REL_MSB                             706
`define DCM_TLAIDTABLEDESC_LKEDCMID_REL_LSB                             700
`define DCM_TLAIDTABLEDESC_LKEDCMID_RESET_VALUE                       7'h64

// macros with short names for field Dcm_TlaIdTableDesc.lkeDcmId
`define DCM_TLIDTBLDSC_LKDCMID_RANGE                                706:700
`define DCM_TLIDTBLDSC_LKDCMID_MSB                                      706
`define DCM_TLIDTBLDSC_LKDCMID_LSB                                      700
`define DCM_TLIDTBLDSC_LKDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_LKDCMID_RESET_VALUE                            7'h64

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.cdeDcmId
`define DCM_TLAIDTABLEDESC_CDEDCMID_RANGE                           713:707
`define DCM_TLAIDTABLEDESC_CDEDCMID_MSB                                 713
`define DCM_TLAIDTABLEDESC_CDEDCMID_LSB                                 707
`define DCM_TLAIDTABLEDESC_CDEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_CDEDCMID_REL_RANGE                       713:707
`define DCM_TLAIDTABLEDESC_CDEDCMID_REL_MSB                             713
`define DCM_TLAIDTABLEDESC_CDEDCMID_REL_LSB                             707
`define DCM_TLAIDTABLEDESC_CDEDCMID_RESET_VALUE                       7'h65

// macros with short names for field Dcm_TlaIdTableDesc.cdeDcmId
`define DCM_TLIDTBLDSC_CDDCMID_RANGE                                713:707
`define DCM_TLIDTBLDSC_CDDCMID_MSB                                      713
`define DCM_TLIDTBLDSC_CDDCMID_LSB                                      707
`define DCM_TLIDTBLDSC_CDDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_CDDCMID_RESET_VALUE                            7'h65

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.nccDcmId
`define DCM_TLAIDTABLEDESC_NCCDCMID_RANGE                           720:714
`define DCM_TLAIDTABLEDESC_NCCDCMID_MSB                                 720
`define DCM_TLAIDTABLEDESC_NCCDCMID_LSB                                 714
`define DCM_TLAIDTABLEDESC_NCCDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NCCDCMID_REL_RANGE                       720:714
`define DCM_TLAIDTABLEDESC_NCCDCMID_REL_MSB                             720
`define DCM_TLAIDTABLEDESC_NCCDCMID_REL_LSB                             714
`define DCM_TLAIDTABLEDESC_NCCDCMID_RESET_VALUE                       7'h66

// macros with short names for field Dcm_TlaIdTableDesc.nccDcmId
`define DCM_TLIDTBLDSC_NCCDCMID_RANGE                               720:714
`define DCM_TLIDTBLDSC_NCCDCMID_MSB                                     720
`define DCM_TLIDTBLDSC_NCCDCMID_LSB                                     714
`define DCM_TLIDTBLDSC_NCCDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_NCCDCMID_RESET_VALUE                           7'h66

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.spqDcmId
`define DCM_TLAIDTABLEDESC_SPQDCMID_RANGE                           727:721
`define DCM_TLAIDTABLEDESC_SPQDCMID_MSB                                 727
`define DCM_TLAIDTABLEDESC_SPQDCMID_LSB                                 721
`define DCM_TLAIDTABLEDESC_SPQDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_SPQDCMID_REL_RANGE                       727:721
`define DCM_TLAIDTABLEDESC_SPQDCMID_REL_MSB                             727
`define DCM_TLAIDTABLEDESC_SPQDCMID_REL_LSB                             721
`define DCM_TLAIDTABLEDESC_SPQDCMID_RESET_VALUE                       7'h67

// macros with short names for field Dcm_TlaIdTableDesc.spqDcmId
`define DCM_TLIDTBLDSC_SPQDCMID_RANGE                               727:721
`define DCM_TLIDTBLDSC_SPQDCMID_MSB                                     727
`define DCM_TLIDTBLDSC_SPQDCMID_LSB                                     721
`define DCM_TLIDTBLDSC_SPQDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_SPQDCMID_RESET_VALUE                           7'h67

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.nmpDcmId
`define DCM_TLAIDTABLEDESC_NMPDCMID_RANGE                           734:728
`define DCM_TLAIDTABLEDESC_NMPDCMID_MSB                                 734
`define DCM_TLAIDTABLEDESC_NMPDCMID_LSB                                 728
`define DCM_TLAIDTABLEDESC_NMPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NMPDCMID_REL_RANGE                       734:728
`define DCM_TLAIDTABLEDESC_NMPDCMID_REL_MSB                             734
`define DCM_TLAIDTABLEDESC_NMPDCMID_REL_LSB                             728
`define DCM_TLAIDTABLEDESC_NMPDCMID_RESET_VALUE                       7'h68

// macros with short names for field Dcm_TlaIdTableDesc.nmpDcmId
`define DCM_TLIDTBLDSC_NMPDCMID_RANGE                               734:728
`define DCM_TLIDTBLDSC_NMPDCMID_MSB                                     734
`define DCM_TLIDTBLDSC_NMPDCMID_LSB                                     728
`define DCM_TLIDTBLDSC_NMPDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_NMPDCMID_RESET_VALUE                           7'h68

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.pxcDcmId
`define DCM_TLAIDTABLEDESC_PXCDCMID_RANGE                           741:735
`define DCM_TLAIDTABLEDESC_PXCDCMID_MSB                                 741
`define DCM_TLAIDTABLEDESC_PXCDCMID_LSB                                 735
`define DCM_TLAIDTABLEDESC_PXCDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_PXCDCMID_REL_RANGE                       741:735
`define DCM_TLAIDTABLEDESC_PXCDCMID_REL_MSB                             741
`define DCM_TLAIDTABLEDESC_PXCDCMID_REL_LSB                             735
`define DCM_TLAIDTABLEDESC_PXCDCMID_RESET_VALUE                       7'h69

// macros with short names for field Dcm_TlaIdTableDesc.pxcDcmId
`define DCM_TLIDTBLDSC_PXCDCMID_RANGE                               741:735
`define DCM_TLIDTBLDSC_PXCDCMID_MSB                                     741
`define DCM_TLIDTBLDSC_PXCDCMID_LSB                                     735
`define DCM_TLIDTBLDSC_PXCDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_PXCDCMID_RESET_VALUE                           7'h69

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.uhdDcmId
`define DCM_TLAIDTABLEDESC_UHDDCMID_RANGE                           748:742
`define DCM_TLAIDTABLEDESC_UHDDCMID_MSB                                 748
`define DCM_TLAIDTABLEDESC_UHDDCMID_LSB                                 742
`define DCM_TLAIDTABLEDESC_UHDDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_UHDDCMID_REL_RANGE                       748:742
`define DCM_TLAIDTABLEDESC_UHDDCMID_REL_MSB                             748
`define DCM_TLAIDTABLEDESC_UHDDCMID_REL_LSB                             742
`define DCM_TLAIDTABLEDESC_UHDDCMID_RESET_VALUE                       7'h6a

// macros with short names for field Dcm_TlaIdTableDesc.uhdDcmId
`define DCM_TLIDTBLDSC_UHDDCMID_RANGE                               748:742
`define DCM_TLIDTBLDSC_UHDDCMID_MSB                                     748
`define DCM_TLIDTBLDSC_UHDDCMID_LSB                                     742
`define DCM_TLIDTBLDSC_UHDDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_UHDDCMID_RESET_VALUE                           7'h6a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ethDcmId
`define DCM_TLAIDTABLEDESC_ETHDCMID_RANGE                           755:749
`define DCM_TLAIDTABLEDESC_ETHDCMID_MSB                                 755
`define DCM_TLAIDTABLEDESC_ETHDCMID_LSB                                 749
`define DCM_TLAIDTABLEDESC_ETHDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_ETHDCMID_REL_RANGE                       755:749
`define DCM_TLAIDTABLEDESC_ETHDCMID_REL_MSB                             755
`define DCM_TLAIDTABLEDESC_ETHDCMID_REL_LSB                             749
`define DCM_TLAIDTABLEDESC_ETHDCMID_RESET_VALUE                       7'h6b

// macros with short names for field Dcm_TlaIdTableDesc.ethDcmId
`define DCM_TLIDTBLDSC_ETHDCMID_RANGE                               755:749
`define DCM_TLIDTBLDSC_ETHDCMID_MSB                                     755
`define DCM_TLIDTBLDSC_ETHDCMID_LSB                                     749
`define DCM_TLIDTBLDSC_ETHDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_ETHDCMID_RESET_VALUE                           7'h6b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ncdDcmId
`define DCM_TLAIDTABLEDESC_NCDDCMID_RANGE                           762:756
`define DCM_TLAIDTABLEDESC_NCDDCMID_MSB                                 762
`define DCM_TLAIDTABLEDESC_NCDDCMID_LSB                                 756
`define DCM_TLAIDTABLEDESC_NCDDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NCDDCMID_REL_RANGE                       762:756
`define DCM_TLAIDTABLEDESC_NCDDCMID_REL_MSB                             762
`define DCM_TLAIDTABLEDESC_NCDDCMID_REL_LSB                             756
`define DCM_TLAIDTABLEDESC_NCDDCMID_RESET_VALUE                       7'h6c

// macros with short names for field Dcm_TlaIdTableDesc.ncdDcmId
`define DCM_TLIDTBLDSC_NCDDCMID_RANGE                               762:756
`define DCM_TLIDTBLDSC_NCDDCMID_MSB                                     762
`define DCM_TLIDTBLDSC_NCDDCMID_LSB                                     756
`define DCM_TLIDTBLDSC_NCDDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_NCDDCMID_RESET_VALUE                           7'h6c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.nspDcmId
`define DCM_TLAIDTABLEDESC_NSPDCMID_RANGE                           769:763
`define DCM_TLAIDTABLEDESC_NSPDCMID_MSB                                 769
`define DCM_TLAIDTABLEDESC_NSPDCMID_LSB                                 763
`define DCM_TLAIDTABLEDESC_NSPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NSPDCMID_REL_RANGE                       769:763
`define DCM_TLAIDTABLEDESC_NSPDCMID_REL_MSB                             769
`define DCM_TLAIDTABLEDESC_NSPDCMID_REL_LSB                             763
`define DCM_TLAIDTABLEDESC_NSPDCMID_RESET_VALUE                       7'h6d

// macros with short names for field Dcm_TlaIdTableDesc.nspDcmId
`define DCM_TLIDTBLDSC_NSPDCMID_RANGE                               769:763
`define DCM_TLIDTBLDSC_NSPDCMID_MSB                                     769
`define DCM_TLIDTBLDSC_NSPDCMID_LSB                                     763
`define DCM_TLIDTBLDSC_NSPDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_NSPDCMID_RESET_VALUE                           7'h6d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.bspDcmId
`define DCM_TLAIDTABLEDESC_BSPDCMID_RANGE                           776:770
`define DCM_TLAIDTABLEDESC_BSPDCMID_MSB                                 776
`define DCM_TLAIDTABLEDESC_BSPDCMID_LSB                                 770
`define DCM_TLAIDTABLEDESC_BSPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_BSPDCMID_REL_RANGE                       776:770
`define DCM_TLAIDTABLEDESC_BSPDCMID_REL_MSB                             776
`define DCM_TLAIDTABLEDESC_BSPDCMID_REL_LSB                             770
`define DCM_TLAIDTABLEDESC_BSPDCMID_RESET_VALUE                       7'h6e

// macros with short names for field Dcm_TlaIdTableDesc.bspDcmId
`define DCM_TLIDTBLDSC_BSPDCMID_RANGE                               776:770
`define DCM_TLIDTBLDSC_BSPDCMID_MSB                                     776
`define DCM_TLIDTBLDSC_BSPDCMID_LSB                                     770
`define DCM_TLIDTBLDSC_BSPDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_BSPDCMID_RESET_VALUE                           7'h6e

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ncaDcmId
`define DCM_TLAIDTABLEDESC_NCADCMID_RANGE                           783:777
`define DCM_TLAIDTABLEDESC_NCADCMID_MSB                                 783
`define DCM_TLAIDTABLEDESC_NCADCMID_LSB                                 777
`define DCM_TLAIDTABLEDESC_NCADCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NCADCMID_REL_RANGE                       783:777
`define DCM_TLAIDTABLEDESC_NCADCMID_REL_MSB                             783
`define DCM_TLAIDTABLEDESC_NCADCMID_REL_LSB                             777
`define DCM_TLAIDTABLEDESC_NCADCMID_RESET_VALUE                       7'h6f

// macros with short names for field Dcm_TlaIdTableDesc.ncaDcmId
`define DCM_TLIDTBLDSC_NCDCMID_RANGE                                783:777
`define DCM_TLIDTBLDSC_NCDCMID_MSB                                      783
`define DCM_TLIDTBLDSC_NCDCMID_LSB                                      777
`define DCM_TLIDTBLDSC_NCDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_NCDCMID_RESET_VALUE                            7'h6f

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.dmcDcmId
`define DCM_TLAIDTABLEDESC_DMCDCMID_RANGE                           790:784
`define DCM_TLAIDTABLEDESC_DMCDCMID_MSB                                 790
`define DCM_TLAIDTABLEDESC_DMCDCMID_LSB                                 784
`define DCM_TLAIDTABLEDESC_DMCDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_DMCDCMID_REL_RANGE                       790:784
`define DCM_TLAIDTABLEDESC_DMCDCMID_REL_MSB                             790
`define DCM_TLAIDTABLEDESC_DMCDCMID_REL_LSB                             784
`define DCM_TLAIDTABLEDESC_DMCDCMID_RESET_VALUE                       7'h70

// macros with short names for field Dcm_TlaIdTableDesc.dmcDcmId
`define DCM_TLIDTBLDSC_DMCDCMID_RANGE                               790:784
`define DCM_TLIDTBLDSC_DMCDCMID_MSB                                     790
`define DCM_TLIDTBLDSC_DMCDCMID_LSB                                     784
`define DCM_TLIDTBLDSC_DMCDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_DMCDCMID_RESET_VALUE                           7'h70

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.nruDcmId
`define DCM_TLAIDTABLEDESC_NRUDCMID_RANGE                           797:791
`define DCM_TLAIDTABLEDESC_NRUDCMID_MSB                                 797
`define DCM_TLAIDTABLEDESC_NRUDCMID_LSB                                 791
`define DCM_TLAIDTABLEDESC_NRUDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NRUDCMID_REL_RANGE                       797:791
`define DCM_TLAIDTABLEDESC_NRUDCMID_REL_MSB                             797
`define DCM_TLAIDTABLEDESC_NRUDCMID_REL_LSB                             791
`define DCM_TLAIDTABLEDESC_NRUDCMID_RESET_VALUE                       7'h71

// macros with short names for field Dcm_TlaIdTableDesc.nruDcmId
`define DCM_TLIDTBLDSC_NRDCMID_RANGE                                797:791
`define DCM_TLIDTBLDSC_NRDCMID_MSB                                      797
`define DCM_TLIDTBLDSC_NRDCMID_LSB                                      791
`define DCM_TLIDTBLDSC_NRDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_NRDCMID_RESET_VALUE                            7'h71

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.xbfDcmId
`define DCM_TLAIDTABLEDESC_XBFDCMID_RANGE                           804:798
`define DCM_TLAIDTABLEDESC_XBFDCMID_MSB                                 804
`define DCM_TLAIDTABLEDESC_XBFDCMID_LSB                                 798
`define DCM_TLAIDTABLEDESC_XBFDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_XBFDCMID_REL_RANGE                       804:798
`define DCM_TLAIDTABLEDESC_XBFDCMID_REL_MSB                             804
`define DCM_TLAIDTABLEDESC_XBFDCMID_REL_LSB                             798
`define DCM_TLAIDTABLEDESC_XBFDCMID_RESET_VALUE                       7'h72

// macros with short names for field Dcm_TlaIdTableDesc.xbfDcmId
`define DCM_TLIDTBLDSC_XBFDCMID_RANGE                               804:798
`define DCM_TLIDTBLDSC_XBFDCMID_MSB                                     804
`define DCM_TLIDTBLDSC_XBFDCMID_LSB                                     798
`define DCM_TLIDTBLDSC_XBFDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_XBFDCMID_RESET_VALUE                           7'h72

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.xbaDcmId
`define DCM_TLAIDTABLEDESC_XBADCMID_RANGE                           811:805
`define DCM_TLAIDTABLEDESC_XBADCMID_MSB                                 811
`define DCM_TLAIDTABLEDESC_XBADCMID_LSB                                 805
`define DCM_TLAIDTABLEDESC_XBADCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_XBADCMID_REL_RANGE                       811:805
`define DCM_TLAIDTABLEDESC_XBADCMID_REL_MSB                             811
`define DCM_TLAIDTABLEDESC_XBADCMID_REL_LSB                             805
`define DCM_TLAIDTABLEDESC_XBADCMID_RESET_VALUE                       7'h73

// macros with short names for field Dcm_TlaIdTableDesc.xbaDcmId
`define DCM_TLIDTBLDSC_XBDCMID_RANGE                                811:805
`define DCM_TLIDTBLDSC_XBDCMID_MSB                                      811
`define DCM_TLIDTBLDSC_XBDCMID_LSB                                      805
`define DCM_TLIDTBLDSC_XBDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_XBDCMID_RESET_VALUE                            7'h73

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.nsiDcmId
`define DCM_TLAIDTABLEDESC_NSIDCMID_RANGE                           818:812
`define DCM_TLAIDTABLEDESC_NSIDCMID_MSB                                 818
`define DCM_TLAIDTABLEDESC_NSIDCMID_LSB                                 812
`define DCM_TLAIDTABLEDESC_NSIDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_NSIDCMID_REL_RANGE                       818:812
`define DCM_TLAIDTABLEDESC_NSIDCMID_REL_MSB                             818
`define DCM_TLAIDTABLEDESC_NSIDCMID_REL_LSB                             812
`define DCM_TLAIDTABLEDESC_NSIDCMID_RESET_VALUE                       7'h74

// macros with short names for field Dcm_TlaIdTableDesc.nsiDcmId
`define DCM_TLIDTBLDSC_NSDCMID_RANGE                                818:812
`define DCM_TLIDTBLDSC_NSDCMID_MSB                                      818
`define DCM_TLIDTBLDSC_NSDCMID_LSB                                      812
`define DCM_TLIDTBLDSC_NSDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_NSDCMID_RESET_VALUE                            7'h74

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.bpiDcmId
`define DCM_TLAIDTABLEDESC_BPIDCMID_RANGE                           825:819
`define DCM_TLAIDTABLEDESC_BPIDCMID_MSB                                 825
`define DCM_TLAIDTABLEDESC_BPIDCMID_LSB                                 819
`define DCM_TLAIDTABLEDESC_BPIDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_BPIDCMID_REL_RANGE                       825:819
`define DCM_TLAIDTABLEDESC_BPIDCMID_REL_MSB                             825
`define DCM_TLAIDTABLEDESC_BPIDCMID_REL_LSB                             819
`define DCM_TLAIDTABLEDESC_BPIDCMID_RESET_VALUE                       7'h75

// macros with short names for field Dcm_TlaIdTableDesc.bpiDcmId
`define DCM_TLIDTBLDSC_BPDCMID_RANGE                                825:819
`define DCM_TLIDTBLDSC_BPDCMID_MSB                                      825
`define DCM_TLIDTBLDSC_BPDCMID_LSB                                      819
`define DCM_TLIDTBLDSC_BPDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_BPDCMID_RESET_VALUE                            7'h75

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.dppDcmId
`define DCM_TLAIDTABLEDESC_DPPDCMID_RANGE                           832:826
`define DCM_TLAIDTABLEDESC_DPPDCMID_MSB                                 832
`define DCM_TLAIDTABLEDESC_DPPDCMID_LSB                                 826
`define DCM_TLAIDTABLEDESC_DPPDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_DPPDCMID_REL_RANGE                       832:826
`define DCM_TLAIDTABLEDESC_DPPDCMID_REL_MSB                             832
`define DCM_TLAIDTABLEDESC_DPPDCMID_REL_LSB                             826
`define DCM_TLAIDTABLEDESC_DPPDCMID_RESET_VALUE                       7'h76

// macros with short names for field Dcm_TlaIdTableDesc.dppDcmId
`define DCM_TLIDTBLDSC_DPPDCMID_RANGE                               832:826
`define DCM_TLIDTBLDSC_DPPDCMID_MSB                                     832
`define DCM_TLIDTBLDSC_DPPDCMID_LSB                                     826
`define DCM_TLIDTBLDSC_DPPDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_DPPDCMID_RESET_VALUE                           7'h76

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.fpxDcmId
`define DCM_TLAIDTABLEDESC_FPXDCMID_RANGE                           839:833
`define DCM_TLAIDTABLEDESC_FPXDCMID_MSB                                 839
`define DCM_TLAIDTABLEDESC_FPXDCMID_LSB                                 833
`define DCM_TLAIDTABLEDESC_FPXDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_FPXDCMID_REL_RANGE                       839:833
`define DCM_TLAIDTABLEDESC_FPXDCMID_REL_MSB                             839
`define DCM_TLAIDTABLEDESC_FPXDCMID_REL_LSB                             833
`define DCM_TLAIDTABLEDESC_FPXDCMID_RESET_VALUE                       7'h77

// macros with short names for field Dcm_TlaIdTableDesc.fpxDcmId
`define DCM_TLIDTBLDSC_FPXDCMID_RANGE                               839:833
`define DCM_TLIDTBLDSC_FPXDCMID_MSB                                     839
`define DCM_TLIDTBLDSC_FPXDCMID_LSB                                     833
`define DCM_TLIDTBLDSC_FPXDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_FPXDCMID_RESET_VALUE                           7'h77

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.hsfDcmId
`define DCM_TLAIDTABLEDESC_HSFDCMID_RANGE                           846:840
`define DCM_TLAIDTABLEDESC_HSFDCMID_MSB                                 846
`define DCM_TLAIDTABLEDESC_HSFDCMID_LSB                                 840
`define DCM_TLAIDTABLEDESC_HSFDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_HSFDCMID_REL_RANGE                       846:840
`define DCM_TLAIDTABLEDESC_HSFDCMID_REL_MSB                             846
`define DCM_TLAIDTABLEDESC_HSFDCMID_REL_LSB                             840
`define DCM_TLAIDTABLEDESC_HSFDCMID_RESET_VALUE                       7'h78

// macros with short names for field Dcm_TlaIdTableDesc.hsfDcmId
`define DCM_TLIDTBLDSC_HSFDCMID_RANGE                               846:840
`define DCM_TLIDTBLDSC_HSFDCMID_MSB                                     846
`define DCM_TLIDTBLDSC_HSFDCMID_LSB                                     840
`define DCM_TLIDTBLDSC_HSFDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_HSFDCMID_RESET_VALUE                           7'h78

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.hsnDcmId
`define DCM_TLAIDTABLEDESC_HSNDCMID_RANGE                           853:847
`define DCM_TLAIDTABLEDESC_HSNDCMID_MSB                                 853
`define DCM_TLAIDTABLEDESC_HSNDCMID_LSB                                 847
`define DCM_TLAIDTABLEDESC_HSNDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_HSNDCMID_REL_RANGE                       853:847
`define DCM_TLAIDTABLEDESC_HSNDCMID_REL_MSB                             853
`define DCM_TLAIDTABLEDESC_HSNDCMID_REL_LSB                             847
`define DCM_TLAIDTABLEDESC_HSNDCMID_RESET_VALUE                       7'h79

// macros with short names for field Dcm_TlaIdTableDesc.hsnDcmId
`define DCM_TLIDTBLDSC_HSNDCMID_RANGE                               853:847
`define DCM_TLIDTBLDSC_HSNDCMID_MSB                                     853
`define DCM_TLIDTBLDSC_HSNDCMID_LSB                                     847
`define DCM_TLIDTBLDSC_HSNDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_HSNDCMID_RESET_VALUE                           7'h79

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.ovfDcmId
`define DCM_TLAIDTABLEDESC_OVFDCMID_RANGE                           860:854
`define DCM_TLAIDTABLEDESC_OVFDCMID_MSB                                 860
`define DCM_TLAIDTABLEDESC_OVFDCMID_LSB                                 854
`define DCM_TLAIDTABLEDESC_OVFDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_OVFDCMID_REL_RANGE                       860:854
`define DCM_TLAIDTABLEDESC_OVFDCMID_REL_MSB                             860
`define DCM_TLAIDTABLEDESC_OVFDCMID_REL_LSB                             854
`define DCM_TLAIDTABLEDESC_OVFDCMID_RESET_VALUE                       7'h7a

// macros with short names for field Dcm_TlaIdTableDesc.ovfDcmId
`define DCM_TLIDTBLDSC_OVFDCMID_RANGE                               860:854
`define DCM_TLIDTBLDSC_OVFDCMID_MSB                                     860
`define DCM_TLIDTBLDSC_OVFDCMID_LSB                                     854
`define DCM_TLIDTBLDSC_OVFDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_OVFDCMID_RESET_VALUE                           7'h7a

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.stcDcmId
`define DCM_TLAIDTABLEDESC_STCDCMID_RANGE                           867:861
`define DCM_TLAIDTABLEDESC_STCDCMID_MSB                                 867
`define DCM_TLAIDTABLEDESC_STCDCMID_LSB                                 861
`define DCM_TLAIDTABLEDESC_STCDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_STCDCMID_REL_RANGE                       867:861
`define DCM_TLAIDTABLEDESC_STCDCMID_REL_MSB                             867
`define DCM_TLAIDTABLEDESC_STCDCMID_REL_LSB                             861
`define DCM_TLAIDTABLEDESC_STCDCMID_RESET_VALUE                       7'h7b

// macros with short names for field Dcm_TlaIdTableDesc.stcDcmId
`define DCM_TLIDTBLDSC_STCDCMID_RANGE                               867:861
`define DCM_TLIDTBLDSC_STCDCMID_MSB                                     867
`define DCM_TLIDTBLDSC_STCDCMID_LSB                                     861
`define DCM_TLIDTBLDSC_STCDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_STCDCMID_RESET_VALUE                           7'h7b

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.stdDcmId
`define DCM_TLAIDTABLEDESC_STDDCMID_RANGE                           874:868
`define DCM_TLAIDTABLEDESC_STDDCMID_MSB                                 874
`define DCM_TLAIDTABLEDESC_STDDCMID_LSB                                 868
`define DCM_TLAIDTABLEDESC_STDDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_STDDCMID_REL_RANGE                       874:868
`define DCM_TLAIDTABLEDESC_STDDCMID_REL_MSB                             874
`define DCM_TLAIDTABLEDESC_STDDCMID_REL_LSB                             868
`define DCM_TLAIDTABLEDESC_STDDCMID_RESET_VALUE                       7'h7c

// macros with short names for field Dcm_TlaIdTableDesc.stdDcmId
`define DCM_TLIDTBLDSC_STDDCMID_RANGE                               874:868
`define DCM_TLIDTBLDSC_STDDCMID_MSB                                     874
`define DCM_TLIDTBLDSC_STDDCMID_LSB                                     868
`define DCM_TLIDTBLDSC_STDDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_STDDCMID_RESET_VALUE                           7'h7c

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.steDcmId
`define DCM_TLAIDTABLEDESC_STEDCMID_RANGE                           881:875
`define DCM_TLAIDTABLEDESC_STEDCMID_MSB                                 881
`define DCM_TLAIDTABLEDESC_STEDCMID_LSB                                 875
`define DCM_TLAIDTABLEDESC_STEDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_STEDCMID_REL_RANGE                       881:875
`define DCM_TLAIDTABLEDESC_STEDCMID_REL_MSB                             881
`define DCM_TLAIDTABLEDESC_STEDCMID_REL_LSB                             875
`define DCM_TLAIDTABLEDESC_STEDCMID_RESET_VALUE                       7'h7d

// macros with short names for field Dcm_TlaIdTableDesc.steDcmId
`define DCM_TLIDTBLDSC_STDCMID_RANGE                                881:875
`define DCM_TLIDTBLDSC_STDCMID_MSB                                      881
`define DCM_TLIDTBLDSC_STDCMID_LSB                                      875
`define DCM_TLIDTBLDSC_STDCMID_WIDTH                                      7
`define DCM_TLIDTBLDSC_STDCMID_RESET_VALUE                            7'h7d

//FieldType - StatusField 
// software : 	 read = true	 write = false	
// hardware : 	 read = true	 write = true	 we = high	
// macros for field Dcm_TlaIdTableDesc.tmqDcmId
`define DCM_TLAIDTABLEDESC_TMQDCMID_RANGE                           888:882
`define DCM_TLAIDTABLEDESC_TMQDCMID_MSB                                 888
`define DCM_TLAIDTABLEDESC_TMQDCMID_LSB                                 882
`define DCM_TLAIDTABLEDESC_TMQDCMID_WIDTH                                 7
`define DCM_TLAIDTABLEDESC_TMQDCMID_REL_RANGE                       888:882
`define DCM_TLAIDTABLEDESC_TMQDCMID_REL_MSB                             888
`define DCM_TLAIDTABLEDESC_TMQDCMID_REL_LSB                             882
`define DCM_TLAIDTABLEDESC_TMQDCMID_RESET_VALUE                       7'h7e

// macros with short names for field Dcm_TlaIdTableDesc.tmqDcmId
`define DCM_TLIDTBLDSC_TMQDCMID_RANGE                               888:882
`define DCM_TLIDTBLDSC_TMQDCMID_MSB                                     888
`define DCM_TLIDTBLDSC_TMQDCMID_LSB                                     882
`define DCM_TLIDTBLDSC_TMQDCMID_WIDTH                                     7
`define DCM_TLIDTBLDSC_TMQDCMID_RESET_VALUE                           7'h7e

//macros for Register - Dcm_TlaIdTableDesc
//Dcm_TlaIdTableDesc is of type DcmTlaIdTableDesc
`define DCM_TLAIDTABLEDESC_REG_NUM                                        1
`define DCM_TLAIDTABLEDESC_REG_ADDR                            32'h00000080
`define DCM_TLAIDTABLEDESC_REG_STRIDE                                   128
`define DCM_TLAIDTABLEDESC_REG_SIZE                                    1024
`define DCM_TLAIDTABLEDESC_REG_FPGA_NUM                                   0
`define DCM_TLAIDTABLEDESC_REG_PHY_SIZE                                 889
`define DCM_TLAIDTABLEDESC_REG_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define DCM_TLAIDTABLEDESC_REG_ADDR_SIZE                                  0
`define DCM_TLAIDTABLEDESC_REG_RESET_VALUE xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx1111110111110111111001111011111101011110011111000111011111101101110101111010011100111110010111000111100001101111110111011011011101100110101111010101101001110100011001111100110110010111001001100011110001011000011100000101111110111101011101101110010110111011010101100110110001010111101011010101011010100101001110100101010001101000010011111001110100110110011001001011100101010010011001000100011110001101000101100010010000111000010100000110000000111111011111001111010111100011101101110100111001011100001101110110110011010101101000110011011001001100010110000010111101011100101101010110001010110101010010100101010000100111010011001001010100100010001101000100100001010000000111110011110001110100111000011011001101000110010011000001011100101100010101001010000100110010010001000100100000001111000111000011010001100000101100010100001001000100000001110000110000010100001000000011000001000000010000000

// macros with short names for register Dcm_TlaIdTableDesc
//Dcm_TlaIdTableDesc is of type DcmTlaIdTableDesc
`define DCM_TLIDTBLDSC_REG_NUM                                            1
`define DCM_TLIDTBLDSC_REG_ADDR                                32'h00000080
`define DCM_TLIDTBLDSC_REG_STRIDE                                       128
`define DCM_TLIDTBLDSC_REG_SIZE                                        1024
`define DCM_TLIDTBLDSC_REG_FPGA_NUM                                       0
`define DCM_TLIDTBLDSC_REG_PHY_SIZE                                     889

`endif // __DCMDESC_VH__
