module ecc_calc (din, eccout);

  parameter ECCDWIDTH = 3;
  parameter ECCWIDTH  = 4;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  generate if (1) begin: inst
    if  (ECCDWIDTH <= 4) 
        ecc_calc_4 ecc_calc (.din(4'b0|din), .eccout(eccout));
    else if  (ECCDWIDTH <= 11)
        ecc_calc_11 ecc_calc (.din(11'b0|din), .eccout(eccout));
    else if  (ECCDWIDTH <= 26)
        ecc_calc_26 ecc_calc (.din(26'b0|din), .eccout(eccout));
    else if  (ECCDWIDTH <= 57)
        ecc_calc_57 ecc_calc (.din(57'b0|din), .eccout(eccout));
    else if  (ECCDWIDTH <= 120)
        ecc_calc_120 ecc_calc (.din(120'b0|din), .eccout(eccout));
    else if  (ECCDWIDTH <= 247)
        ecc_calc_247 ecc_calc (.din(247'b0|din), .eccout(eccout));
    else if  (ECCDWIDTH <= 502)
        ecc_calc_502 ecc_calc (.din(502'b0|din), .eccout(eccout));
  end
  endgenerate

endmodule

module ecc_calc_4 (din, eccout);

  localparam ECCDWIDTH = 4;
  localparam ECCWIDTH  = 4;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  wire [ECCDWIDTH-1:0]   ecchmatrix [0:ECCWIDTH-1];

 assign eccout[3] = ^(ecchmatrix[3]&din);
 assign eccout[2] = ^(ecchmatrix[2]&din);
 assign eccout[1] = ^(ecchmatrix[1]&din);
 assign eccout[0] = ^(ecchmatrix[0]&din);
// assign ready = 1'b1;

// Generate the H Matrix in Perl

// Initialize the hmatrix array
   assign ecchmatrix[0][0] = 1;
   assign ecchmatrix[1][0] = 1;
   assign ecchmatrix[2][0] = 1;
   assign ecchmatrix[3][0] = 0;
   assign ecchmatrix[0][1] = 1;
   assign ecchmatrix[1][1] = 1;
   assign ecchmatrix[2][1] = 0;
   assign ecchmatrix[3][1] = 1;
   assign ecchmatrix[0][2] = 1;
   assign ecchmatrix[1][2] = 0;
   assign ecchmatrix[2][2] = 1;
   assign ecchmatrix[3][2] = 1;
   assign ecchmatrix[0][3] = 0;
   assign ecchmatrix[1][3] = 1;
   assign ecchmatrix[2][3] = 1;
   assign ecchmatrix[3][3] = 1;
endmodule

module ecc_calc_11 (din, eccout);

  localparam ECCDWIDTH = 11;
  localparam ECCWIDTH  = 5;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  wire [ECCDWIDTH-1:0]   ecchmatrix [0:ECCWIDTH-1];

 assign eccout[4] = ^(ecchmatrix[4]&din);
 assign eccout[3] = ^(ecchmatrix[3]&din);
 assign eccout[2] = ^(ecchmatrix[2]&din);
 assign eccout[1] = ^(ecchmatrix[1]&din);
 assign eccout[0] = ^(ecchmatrix[0]&din);
// assign ready = 1'b1;

// Generate the H Matrix in Perl

// Initialize the hmatrix array
   assign ecchmatrix[0][0] = 1;
   assign ecchmatrix[1][0] = 1;
   assign ecchmatrix[2][0] = 1;
   assign ecchmatrix[3][0] = 0;
   assign ecchmatrix[4][0] = 0;
   assign ecchmatrix[0][1] = 1;
   assign ecchmatrix[1][1] = 1;
   assign ecchmatrix[2][1] = 0;
   assign ecchmatrix[3][1] = 1;
   assign ecchmatrix[4][1] = 0;
   assign ecchmatrix[0][2] = 1;
   assign ecchmatrix[1][2] = 1;
   assign ecchmatrix[2][2] = 0;
   assign ecchmatrix[3][2] = 0;
   assign ecchmatrix[4][2] = 1;
   assign ecchmatrix[0][3] = 1;
   assign ecchmatrix[1][3] = 0;
   assign ecchmatrix[2][3] = 1;
   assign ecchmatrix[3][3] = 1;
   assign ecchmatrix[4][3] = 0;
   assign ecchmatrix[0][4] = 1;
   assign ecchmatrix[1][4] = 0;
   assign ecchmatrix[2][4] = 1;
   assign ecchmatrix[3][4] = 0;
   assign ecchmatrix[4][4] = 1;
   assign ecchmatrix[0][5] = 1;
   assign ecchmatrix[1][5] = 0;
   assign ecchmatrix[2][5] = 0;
   assign ecchmatrix[3][5] = 1;
   assign ecchmatrix[4][5] = 1;
   assign ecchmatrix[0][6] = 0;
   assign ecchmatrix[1][6] = 1;
   assign ecchmatrix[2][6] = 1;
   assign ecchmatrix[3][6] = 1;
   assign ecchmatrix[4][6] = 0;
   assign ecchmatrix[0][7] = 0;
   assign ecchmatrix[1][7] = 1;
   assign ecchmatrix[2][7] = 1;
   assign ecchmatrix[3][7] = 0;
   assign ecchmatrix[4][7] = 1;
   assign ecchmatrix[0][8] = 0;
   assign ecchmatrix[1][8] = 1;
   assign ecchmatrix[2][8] = 0;
   assign ecchmatrix[3][8] = 1;
   assign ecchmatrix[4][8] = 1;
   assign ecchmatrix[0][9] = 0;
   assign ecchmatrix[1][9] = 0;
   assign ecchmatrix[2][9] = 1;
   assign ecchmatrix[3][9] = 1;
   assign ecchmatrix[4][9] = 1;
   assign ecchmatrix[0][10] = 1;
   assign ecchmatrix[1][10] = 1;
   assign ecchmatrix[2][10] = 1;
   assign ecchmatrix[3][10] = 1;
   assign ecchmatrix[4][10] = 1;
endmodule

module ecc_calc_26 (din, eccout);

  localparam ECCDWIDTH = 26;
  localparam ECCWIDTH  = 6;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  wire [ECCDWIDTH-1:0]   ecchmatrix [0:ECCWIDTH-1];

 assign eccout[5] = ^(ecchmatrix[5]&din);
 assign eccout[4] = ^(ecchmatrix[4]&din);
 assign eccout[3] = ^(ecchmatrix[3]&din);
 assign eccout[2] = ^(ecchmatrix[2]&din);
 assign eccout[1] = ^(ecchmatrix[1]&din);
 assign eccout[0] = ^(ecchmatrix[0]&din);
// assign ready = 1'b1;

// Generate the H Matrix in Perl

// Initialize the hmatrix array
   assign ecchmatrix[0][0] = 1;
   assign ecchmatrix[1][0] = 1;
   assign ecchmatrix[2][0] = 1;
   assign ecchmatrix[3][0] = 0;
   assign ecchmatrix[4][0] = 0;
   assign ecchmatrix[5][0] = 0;
   assign ecchmatrix[0][1] = 1;
   assign ecchmatrix[1][1] = 1;
   assign ecchmatrix[2][1] = 0;
   assign ecchmatrix[3][1] = 1;
   assign ecchmatrix[4][1] = 0;
   assign ecchmatrix[5][1] = 0;
   assign ecchmatrix[0][2] = 1;
   assign ecchmatrix[1][2] = 1;
   assign ecchmatrix[2][2] = 0;
   assign ecchmatrix[3][2] = 0;
   assign ecchmatrix[4][2] = 1;
   assign ecchmatrix[5][2] = 0;
   assign ecchmatrix[0][3] = 1;
   assign ecchmatrix[1][3] = 1;
   assign ecchmatrix[2][3] = 0;
   assign ecchmatrix[3][3] = 0;
   assign ecchmatrix[4][3] = 0;
   assign ecchmatrix[5][3] = 1;
   assign ecchmatrix[0][4] = 1;
   assign ecchmatrix[1][4] = 0;
   assign ecchmatrix[2][4] = 1;
   assign ecchmatrix[3][4] = 1;
   assign ecchmatrix[4][4] = 0;
   assign ecchmatrix[5][4] = 0;
   assign ecchmatrix[0][5] = 1;
   assign ecchmatrix[1][5] = 0;
   assign ecchmatrix[2][5] = 1;
   assign ecchmatrix[3][5] = 0;
   assign ecchmatrix[4][5] = 1;
   assign ecchmatrix[5][5] = 0;
   assign ecchmatrix[0][6] = 1;
   assign ecchmatrix[1][6] = 0;
   assign ecchmatrix[2][6] = 1;
   assign ecchmatrix[3][6] = 0;
   assign ecchmatrix[4][6] = 0;
   assign ecchmatrix[5][6] = 1;
   assign ecchmatrix[0][7] = 1;
   assign ecchmatrix[1][7] = 0;
   assign ecchmatrix[2][7] = 0;
   assign ecchmatrix[3][7] = 1;
   assign ecchmatrix[4][7] = 1;
   assign ecchmatrix[5][7] = 0;
   assign ecchmatrix[0][8] = 1;
   assign ecchmatrix[1][8] = 0;
   assign ecchmatrix[2][8] = 0;
   assign ecchmatrix[3][8] = 1;
   assign ecchmatrix[4][8] = 0;
   assign ecchmatrix[5][8] = 1;
   assign ecchmatrix[0][9] = 1;
   assign ecchmatrix[1][9] = 0;
   assign ecchmatrix[2][9] = 0;
   assign ecchmatrix[3][9] = 0;
   assign ecchmatrix[4][9] = 1;
   assign ecchmatrix[5][9] = 1;
   assign ecchmatrix[0][10] = 0;
   assign ecchmatrix[1][10] = 1;
   assign ecchmatrix[2][10] = 1;
   assign ecchmatrix[3][10] = 1;
   assign ecchmatrix[4][10] = 0;
   assign ecchmatrix[5][10] = 0;
   assign ecchmatrix[0][11] = 0;
   assign ecchmatrix[1][11] = 1;
   assign ecchmatrix[2][11] = 1;
   assign ecchmatrix[3][11] = 0;
   assign ecchmatrix[4][11] = 1;
   assign ecchmatrix[5][11] = 0;
   assign ecchmatrix[0][12] = 0;
   assign ecchmatrix[1][12] = 1;
   assign ecchmatrix[2][12] = 1;
   assign ecchmatrix[3][12] = 0;
   assign ecchmatrix[4][12] = 0;
   assign ecchmatrix[5][12] = 1;
   assign ecchmatrix[0][13] = 0;
   assign ecchmatrix[1][13] = 1;
   assign ecchmatrix[2][13] = 0;
   assign ecchmatrix[3][13] = 1;
   assign ecchmatrix[4][13] = 1;
   assign ecchmatrix[5][13] = 0;
   assign ecchmatrix[0][14] = 0;
   assign ecchmatrix[1][14] = 1;
   assign ecchmatrix[2][14] = 0;
   assign ecchmatrix[3][14] = 1;
   assign ecchmatrix[4][14] = 0;
   assign ecchmatrix[5][14] = 1;
   assign ecchmatrix[0][15] = 0;
   assign ecchmatrix[1][15] = 1;
   assign ecchmatrix[2][15] = 0;
   assign ecchmatrix[3][15] = 0;
   assign ecchmatrix[4][15] = 1;
   assign ecchmatrix[5][15] = 1;
   assign ecchmatrix[0][16] = 0;
   assign ecchmatrix[1][16] = 0;
   assign ecchmatrix[2][16] = 1;
   assign ecchmatrix[3][16] = 1;
   assign ecchmatrix[4][16] = 1;
   assign ecchmatrix[5][16] = 0;
   assign ecchmatrix[0][17] = 0;
   assign ecchmatrix[1][17] = 0;
   assign ecchmatrix[2][17] = 1;
   assign ecchmatrix[3][17] = 1;
   assign ecchmatrix[4][17] = 0;
   assign ecchmatrix[5][17] = 1;
   assign ecchmatrix[0][18] = 0;
   assign ecchmatrix[1][18] = 0;
   assign ecchmatrix[2][18] = 1;
   assign ecchmatrix[3][18] = 0;
   assign ecchmatrix[4][18] = 1;
   assign ecchmatrix[5][18] = 1;
   assign ecchmatrix[0][19] = 0;
   assign ecchmatrix[1][19] = 0;
   assign ecchmatrix[2][19] = 0;
   assign ecchmatrix[3][19] = 1;
   assign ecchmatrix[4][19] = 1;
   assign ecchmatrix[5][19] = 1;
   assign ecchmatrix[0][20] = 1;
   assign ecchmatrix[1][20] = 1;
   assign ecchmatrix[2][20] = 1;
   assign ecchmatrix[3][20] = 1;
   assign ecchmatrix[4][20] = 1;
   assign ecchmatrix[5][20] = 0;
   assign ecchmatrix[0][21] = 1;
   assign ecchmatrix[1][21] = 1;
   assign ecchmatrix[2][21] = 1;
   assign ecchmatrix[3][21] = 1;
   assign ecchmatrix[4][21] = 0;
   assign ecchmatrix[5][21] = 1;
   assign ecchmatrix[0][22] = 1;
   assign ecchmatrix[1][22] = 1;
   assign ecchmatrix[2][22] = 1;
   assign ecchmatrix[3][22] = 0;
   assign ecchmatrix[4][22] = 1;
   assign ecchmatrix[5][22] = 1;
   assign ecchmatrix[0][23] = 1;
   assign ecchmatrix[1][23] = 1;
   assign ecchmatrix[2][23] = 0;
   assign ecchmatrix[3][23] = 1;
   assign ecchmatrix[4][23] = 1;
   assign ecchmatrix[5][23] = 1;
   assign ecchmatrix[0][24] = 1;
   assign ecchmatrix[1][24] = 0;
   assign ecchmatrix[2][24] = 1;
   assign ecchmatrix[3][24] = 1;
   assign ecchmatrix[4][24] = 1;
   assign ecchmatrix[5][24] = 1;
   assign ecchmatrix[0][25] = 0;
   assign ecchmatrix[1][25] = 1;
   assign ecchmatrix[2][25] = 1;
   assign ecchmatrix[3][25] = 1;
   assign ecchmatrix[4][25] = 1;
   assign ecchmatrix[5][25] = 1;
endmodule

module ecc_calc_57 (din, eccout);

  localparam ECCDWIDTH = 57;
  localparam ECCWIDTH  = 7;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  wire [ECCDWIDTH-1:0]   ecchmatrix [0:ECCWIDTH-1];

 assign eccout[6] = ^(ecchmatrix[6]&din);
 assign eccout[5] = ^(ecchmatrix[5]&din);
 assign eccout[4] = ^(ecchmatrix[4]&din);
 assign eccout[3] = ^(ecchmatrix[3]&din);
 assign eccout[2] = ^(ecchmatrix[2]&din);
 assign eccout[1] = ^(ecchmatrix[1]&din);
 assign eccout[0] = ^(ecchmatrix[0]&din);
// assign ready = 1'b1;

// Generate the H Matrix in Perl

// Initialize the hmatrix array
   assign ecchmatrix[0][0] = 1;
   assign ecchmatrix[1][0] = 1;
   assign ecchmatrix[2][0] = 1;
   assign ecchmatrix[3][0] = 0;
   assign ecchmatrix[4][0] = 0;
   assign ecchmatrix[5][0] = 0;
   assign ecchmatrix[6][0] = 0;
   assign ecchmatrix[0][1] = 1;
   assign ecchmatrix[1][1] = 1;
   assign ecchmatrix[2][1] = 0;
   assign ecchmatrix[3][1] = 1;
   assign ecchmatrix[4][1] = 0;
   assign ecchmatrix[5][1] = 0;
   assign ecchmatrix[6][1] = 0;
   assign ecchmatrix[0][2] = 1;
   assign ecchmatrix[1][2] = 1;
   assign ecchmatrix[2][2] = 0;
   assign ecchmatrix[3][2] = 0;
   assign ecchmatrix[4][2] = 1;
   assign ecchmatrix[5][2] = 0;
   assign ecchmatrix[6][2] = 0;
   assign ecchmatrix[0][3] = 1;
   assign ecchmatrix[1][3] = 1;
   assign ecchmatrix[2][3] = 0;
   assign ecchmatrix[3][3] = 0;
   assign ecchmatrix[4][3] = 0;
   assign ecchmatrix[5][3] = 1;
   assign ecchmatrix[6][3] = 0;
   assign ecchmatrix[0][4] = 1;
   assign ecchmatrix[1][4] = 1;
   assign ecchmatrix[2][4] = 0;
   assign ecchmatrix[3][4] = 0;
   assign ecchmatrix[4][4] = 0;
   assign ecchmatrix[5][4] = 0;
   assign ecchmatrix[6][4] = 1;
   assign ecchmatrix[0][5] = 1;
   assign ecchmatrix[1][5] = 0;
   assign ecchmatrix[2][5] = 1;
   assign ecchmatrix[3][5] = 1;
   assign ecchmatrix[4][5] = 0;
   assign ecchmatrix[5][5] = 0;
   assign ecchmatrix[6][5] = 0;
   assign ecchmatrix[0][6] = 1;
   assign ecchmatrix[1][6] = 0;
   assign ecchmatrix[2][6] = 1;
   assign ecchmatrix[3][6] = 0;
   assign ecchmatrix[4][6] = 1;
   assign ecchmatrix[5][6] = 0;
   assign ecchmatrix[6][6] = 0;
   assign ecchmatrix[0][7] = 1;
   assign ecchmatrix[1][7] = 0;
   assign ecchmatrix[2][7] = 1;
   assign ecchmatrix[3][7] = 0;
   assign ecchmatrix[4][7] = 0;
   assign ecchmatrix[5][7] = 1;
   assign ecchmatrix[6][7] = 0;
   assign ecchmatrix[0][8] = 1;
   assign ecchmatrix[1][8] = 0;
   assign ecchmatrix[2][8] = 1;
   assign ecchmatrix[3][8] = 0;
   assign ecchmatrix[4][8] = 0;
   assign ecchmatrix[5][8] = 0;
   assign ecchmatrix[6][8] = 1;
   assign ecchmatrix[0][9] = 1;
   assign ecchmatrix[1][9] = 0;
   assign ecchmatrix[2][9] = 0;
   assign ecchmatrix[3][9] = 1;
   assign ecchmatrix[4][9] = 1;
   assign ecchmatrix[5][9] = 0;
   assign ecchmatrix[6][9] = 0;
   assign ecchmatrix[0][10] = 1;
   assign ecchmatrix[1][10] = 0;
   assign ecchmatrix[2][10] = 0;
   assign ecchmatrix[3][10] = 1;
   assign ecchmatrix[4][10] = 0;
   assign ecchmatrix[5][10] = 1;
   assign ecchmatrix[6][10] = 0;
   assign ecchmatrix[0][11] = 1;
   assign ecchmatrix[1][11] = 0;
   assign ecchmatrix[2][11] = 0;
   assign ecchmatrix[3][11] = 1;
   assign ecchmatrix[4][11] = 0;
   assign ecchmatrix[5][11] = 0;
   assign ecchmatrix[6][11] = 1;
   assign ecchmatrix[0][12] = 1;
   assign ecchmatrix[1][12] = 0;
   assign ecchmatrix[2][12] = 0;
   assign ecchmatrix[3][12] = 0;
   assign ecchmatrix[4][12] = 1;
   assign ecchmatrix[5][12] = 1;
   assign ecchmatrix[6][12] = 0;
   assign ecchmatrix[0][13] = 1;
   assign ecchmatrix[1][13] = 0;
   assign ecchmatrix[2][13] = 0;
   assign ecchmatrix[3][13] = 0;
   assign ecchmatrix[4][13] = 1;
   assign ecchmatrix[5][13] = 0;
   assign ecchmatrix[6][13] = 1;
   assign ecchmatrix[0][14] = 1;
   assign ecchmatrix[1][14] = 0;
   assign ecchmatrix[2][14] = 0;
   assign ecchmatrix[3][14] = 0;
   assign ecchmatrix[4][14] = 0;
   assign ecchmatrix[5][14] = 1;
   assign ecchmatrix[6][14] = 1;
   assign ecchmatrix[0][15] = 0;
   assign ecchmatrix[1][15] = 1;
   assign ecchmatrix[2][15] = 1;
   assign ecchmatrix[3][15] = 1;
   assign ecchmatrix[4][15] = 0;
   assign ecchmatrix[5][15] = 0;
   assign ecchmatrix[6][15] = 0;
   assign ecchmatrix[0][16] = 0;
   assign ecchmatrix[1][16] = 1;
   assign ecchmatrix[2][16] = 1;
   assign ecchmatrix[3][16] = 0;
   assign ecchmatrix[4][16] = 1;
   assign ecchmatrix[5][16] = 0;
   assign ecchmatrix[6][16] = 0;
   assign ecchmatrix[0][17] = 0;
   assign ecchmatrix[1][17] = 1;
   assign ecchmatrix[2][17] = 1;
   assign ecchmatrix[3][17] = 0;
   assign ecchmatrix[4][17] = 0;
   assign ecchmatrix[5][17] = 1;
   assign ecchmatrix[6][17] = 0;
   assign ecchmatrix[0][18] = 0;
   assign ecchmatrix[1][18] = 1;
   assign ecchmatrix[2][18] = 1;
   assign ecchmatrix[3][18] = 0;
   assign ecchmatrix[4][18] = 0;
   assign ecchmatrix[5][18] = 0;
   assign ecchmatrix[6][18] = 1;
   assign ecchmatrix[0][19] = 0;
   assign ecchmatrix[1][19] = 1;
   assign ecchmatrix[2][19] = 0;
   assign ecchmatrix[3][19] = 1;
   assign ecchmatrix[4][19] = 1;
   assign ecchmatrix[5][19] = 0;
   assign ecchmatrix[6][19] = 0;
   assign ecchmatrix[0][20] = 0;
   assign ecchmatrix[1][20] = 1;
   assign ecchmatrix[2][20] = 0;
   assign ecchmatrix[3][20] = 1;
   assign ecchmatrix[4][20] = 0;
   assign ecchmatrix[5][20] = 1;
   assign ecchmatrix[6][20] = 0;
   assign ecchmatrix[0][21] = 0;
   assign ecchmatrix[1][21] = 1;
   assign ecchmatrix[2][21] = 0;
   assign ecchmatrix[3][21] = 1;
   assign ecchmatrix[4][21] = 0;
   assign ecchmatrix[5][21] = 0;
   assign ecchmatrix[6][21] = 1;
   assign ecchmatrix[0][22] = 0;
   assign ecchmatrix[1][22] = 1;
   assign ecchmatrix[2][22] = 0;
   assign ecchmatrix[3][22] = 0;
   assign ecchmatrix[4][22] = 1;
   assign ecchmatrix[5][22] = 1;
   assign ecchmatrix[6][22] = 0;
   assign ecchmatrix[0][23] = 0;
   assign ecchmatrix[1][23] = 1;
   assign ecchmatrix[2][23] = 0;
   assign ecchmatrix[3][23] = 0;
   assign ecchmatrix[4][23] = 1;
   assign ecchmatrix[5][23] = 0;
   assign ecchmatrix[6][23] = 1;
   assign ecchmatrix[0][24] = 0;
   assign ecchmatrix[1][24] = 1;
   assign ecchmatrix[2][24] = 0;
   assign ecchmatrix[3][24] = 0;
   assign ecchmatrix[4][24] = 0;
   assign ecchmatrix[5][24] = 1;
   assign ecchmatrix[6][24] = 1;
   assign ecchmatrix[0][25] = 0;
   assign ecchmatrix[1][25] = 0;
   assign ecchmatrix[2][25] = 1;
   assign ecchmatrix[3][25] = 1;
   assign ecchmatrix[4][25] = 1;
   assign ecchmatrix[5][25] = 0;
   assign ecchmatrix[6][25] = 0;
   assign ecchmatrix[0][26] = 0;
   assign ecchmatrix[1][26] = 0;
   assign ecchmatrix[2][26] = 1;
   assign ecchmatrix[3][26] = 1;
   assign ecchmatrix[4][26] = 0;
   assign ecchmatrix[5][26] = 1;
   assign ecchmatrix[6][26] = 0;
   assign ecchmatrix[0][27] = 0;
   assign ecchmatrix[1][27] = 0;
   assign ecchmatrix[2][27] = 1;
   assign ecchmatrix[3][27] = 1;
   assign ecchmatrix[4][27] = 0;
   assign ecchmatrix[5][27] = 0;
   assign ecchmatrix[6][27] = 1;
   assign ecchmatrix[0][28] = 0;
   assign ecchmatrix[1][28] = 0;
   assign ecchmatrix[2][28] = 1;
   assign ecchmatrix[3][28] = 0;
   assign ecchmatrix[4][28] = 1;
   assign ecchmatrix[5][28] = 1;
   assign ecchmatrix[6][28] = 0;
   assign ecchmatrix[0][29] = 0;
   assign ecchmatrix[1][29] = 0;
   assign ecchmatrix[2][29] = 1;
   assign ecchmatrix[3][29] = 0;
   assign ecchmatrix[4][29] = 1;
   assign ecchmatrix[5][29] = 0;
   assign ecchmatrix[6][29] = 1;
   assign ecchmatrix[0][30] = 0;
   assign ecchmatrix[1][30] = 0;
   assign ecchmatrix[2][30] = 1;
   assign ecchmatrix[3][30] = 0;
   assign ecchmatrix[4][30] = 0;
   assign ecchmatrix[5][30] = 1;
   assign ecchmatrix[6][30] = 1;
   assign ecchmatrix[0][31] = 0;
   assign ecchmatrix[1][31] = 0;
   assign ecchmatrix[2][31] = 0;
   assign ecchmatrix[3][31] = 1;
   assign ecchmatrix[4][31] = 1;
   assign ecchmatrix[5][31] = 1;
   assign ecchmatrix[6][31] = 0;
   assign ecchmatrix[0][32] = 0;
   assign ecchmatrix[1][32] = 0;
   assign ecchmatrix[2][32] = 0;
   assign ecchmatrix[3][32] = 1;
   assign ecchmatrix[4][32] = 1;
   assign ecchmatrix[5][32] = 0;
   assign ecchmatrix[6][32] = 1;
   assign ecchmatrix[0][33] = 0;
   assign ecchmatrix[1][33] = 0;
   assign ecchmatrix[2][33] = 0;
   assign ecchmatrix[3][33] = 1;
   assign ecchmatrix[4][33] = 0;
   assign ecchmatrix[5][33] = 1;
   assign ecchmatrix[6][33] = 1;
   assign ecchmatrix[0][34] = 0;
   assign ecchmatrix[1][34] = 0;
   assign ecchmatrix[2][34] = 0;
   assign ecchmatrix[3][34] = 0;
   assign ecchmatrix[4][34] = 1;
   assign ecchmatrix[5][34] = 1;
   assign ecchmatrix[6][34] = 1;
   assign ecchmatrix[0][35] = 1;
   assign ecchmatrix[1][35] = 1;
   assign ecchmatrix[2][35] = 1;
   assign ecchmatrix[3][35] = 1;
   assign ecchmatrix[4][35] = 1;
   assign ecchmatrix[5][35] = 0;
   assign ecchmatrix[6][35] = 0;
   assign ecchmatrix[0][36] = 1;
   assign ecchmatrix[1][36] = 1;
   assign ecchmatrix[2][36] = 1;
   assign ecchmatrix[3][36] = 1;
   assign ecchmatrix[4][36] = 0;
   assign ecchmatrix[5][36] = 1;
   assign ecchmatrix[6][36] = 0;
   assign ecchmatrix[0][37] = 1;
   assign ecchmatrix[1][37] = 1;
   assign ecchmatrix[2][37] = 1;
   assign ecchmatrix[3][37] = 1;
   assign ecchmatrix[4][37] = 0;
   assign ecchmatrix[5][37] = 0;
   assign ecchmatrix[6][37] = 1;
   assign ecchmatrix[0][38] = 1;
   assign ecchmatrix[1][38] = 1;
   assign ecchmatrix[2][38] = 1;
   assign ecchmatrix[3][38] = 0;
   assign ecchmatrix[4][38] = 1;
   assign ecchmatrix[5][38] = 1;
   assign ecchmatrix[6][38] = 0;
   assign ecchmatrix[0][39] = 1;
   assign ecchmatrix[1][39] = 1;
   assign ecchmatrix[2][39] = 1;
   assign ecchmatrix[3][39] = 0;
   assign ecchmatrix[4][39] = 1;
   assign ecchmatrix[5][39] = 0;
   assign ecchmatrix[6][39] = 1;
   assign ecchmatrix[0][40] = 1;
   assign ecchmatrix[1][40] = 1;
   assign ecchmatrix[2][40] = 1;
   assign ecchmatrix[3][40] = 0;
   assign ecchmatrix[4][40] = 0;
   assign ecchmatrix[5][40] = 1;
   assign ecchmatrix[6][40] = 1;
   assign ecchmatrix[0][41] = 1;
   assign ecchmatrix[1][41] = 1;
   assign ecchmatrix[2][41] = 0;
   assign ecchmatrix[3][41] = 1;
   assign ecchmatrix[4][41] = 1;
   assign ecchmatrix[5][41] = 1;
   assign ecchmatrix[6][41] = 0;
   assign ecchmatrix[0][42] = 1;
   assign ecchmatrix[1][42] = 1;
   assign ecchmatrix[2][42] = 0;
   assign ecchmatrix[3][42] = 1;
   assign ecchmatrix[4][42] = 1;
   assign ecchmatrix[5][42] = 0;
   assign ecchmatrix[6][42] = 1;
   assign ecchmatrix[0][43] = 1;
   assign ecchmatrix[1][43] = 1;
   assign ecchmatrix[2][43] = 0;
   assign ecchmatrix[3][43] = 1;
   assign ecchmatrix[4][43] = 0;
   assign ecchmatrix[5][43] = 1;
   assign ecchmatrix[6][43] = 1;
   assign ecchmatrix[0][44] = 1;
   assign ecchmatrix[1][44] = 1;
   assign ecchmatrix[2][44] = 0;
   assign ecchmatrix[3][44] = 0;
   assign ecchmatrix[4][44] = 1;
   assign ecchmatrix[5][44] = 1;
   assign ecchmatrix[6][44] = 1;
   assign ecchmatrix[0][45] = 1;
   assign ecchmatrix[1][45] = 0;
   assign ecchmatrix[2][45] = 1;
   assign ecchmatrix[3][45] = 1;
   assign ecchmatrix[4][45] = 1;
   assign ecchmatrix[5][45] = 1;
   assign ecchmatrix[6][45] = 0;
   assign ecchmatrix[0][46] = 1;
   assign ecchmatrix[1][46] = 0;
   assign ecchmatrix[2][46] = 1;
   assign ecchmatrix[3][46] = 1;
   assign ecchmatrix[4][46] = 1;
   assign ecchmatrix[5][46] = 0;
   assign ecchmatrix[6][46] = 1;
   assign ecchmatrix[0][47] = 1;
   assign ecchmatrix[1][47] = 0;
   assign ecchmatrix[2][47] = 1;
   assign ecchmatrix[3][47] = 1;
   assign ecchmatrix[4][47] = 0;
   assign ecchmatrix[5][47] = 1;
   assign ecchmatrix[6][47] = 1;
   assign ecchmatrix[0][48] = 1;
   assign ecchmatrix[1][48] = 0;
   assign ecchmatrix[2][48] = 1;
   assign ecchmatrix[3][48] = 0;
   assign ecchmatrix[4][48] = 1;
   assign ecchmatrix[5][48] = 1;
   assign ecchmatrix[6][48] = 1;
   assign ecchmatrix[0][49] = 1;
   assign ecchmatrix[1][49] = 0;
   assign ecchmatrix[2][49] = 0;
   assign ecchmatrix[3][49] = 1;
   assign ecchmatrix[4][49] = 1;
   assign ecchmatrix[5][49] = 1;
   assign ecchmatrix[6][49] = 1;
   assign ecchmatrix[0][50] = 0;
   assign ecchmatrix[1][50] = 1;
   assign ecchmatrix[2][50] = 1;
   assign ecchmatrix[3][50] = 1;
   assign ecchmatrix[4][50] = 1;
   assign ecchmatrix[5][50] = 1;
   assign ecchmatrix[6][50] = 0;
   assign ecchmatrix[0][51] = 0;
   assign ecchmatrix[1][51] = 1;
   assign ecchmatrix[2][51] = 1;
   assign ecchmatrix[3][51] = 1;
   assign ecchmatrix[4][51] = 1;
   assign ecchmatrix[5][51] = 0;
   assign ecchmatrix[6][51] = 1;
   assign ecchmatrix[0][52] = 0;
   assign ecchmatrix[1][52] = 1;
   assign ecchmatrix[2][52] = 1;
   assign ecchmatrix[3][52] = 1;
   assign ecchmatrix[4][52] = 0;
   assign ecchmatrix[5][52] = 1;
   assign ecchmatrix[6][52] = 1;
   assign ecchmatrix[0][53] = 0;
   assign ecchmatrix[1][53] = 1;
   assign ecchmatrix[2][53] = 1;
   assign ecchmatrix[3][53] = 0;
   assign ecchmatrix[4][53] = 1;
   assign ecchmatrix[5][53] = 1;
   assign ecchmatrix[6][53] = 1;
   assign ecchmatrix[0][54] = 0;
   assign ecchmatrix[1][54] = 1;
   assign ecchmatrix[2][54] = 0;
   assign ecchmatrix[3][54] = 1;
   assign ecchmatrix[4][54] = 1;
   assign ecchmatrix[5][54] = 1;
   assign ecchmatrix[6][54] = 1;
   assign ecchmatrix[0][55] = 0;
   assign ecchmatrix[1][55] = 0;
   assign ecchmatrix[2][55] = 1;
   assign ecchmatrix[3][55] = 1;
   assign ecchmatrix[4][55] = 1;
   assign ecchmatrix[5][55] = 1;
   assign ecchmatrix[6][55] = 1;
   assign ecchmatrix[0][56] = 1;
   assign ecchmatrix[1][56] = 1;
   assign ecchmatrix[2][56] = 1;
   assign ecchmatrix[3][56] = 1;
   assign ecchmatrix[4][56] = 1;
   assign ecchmatrix[5][56] = 1;
   assign ecchmatrix[6][56] = 1;
endmodule

module ecc_calc_120 (din, eccout);

  localparam ECCDWIDTH = 120;
  localparam ECCWIDTH  = 8;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  wire [ECCDWIDTH-1:0]   ecchmatrix [0:ECCWIDTH-1];

 assign eccout[7] = ^(ecchmatrix[7]&din);
 assign eccout[6] = ^(ecchmatrix[6]&din);
 assign eccout[5] = ^(ecchmatrix[5]&din);
 assign eccout[4] = ^(ecchmatrix[4]&din);
 assign eccout[3] = ^(ecchmatrix[3]&din);
 assign eccout[2] = ^(ecchmatrix[2]&din);
 assign eccout[1] = ^(ecchmatrix[1]&din);
 assign eccout[0] = ^(ecchmatrix[0]&din);
// assign ready = 1'b1;

// Generate the H Matrix in Perl

// Initialize the hmatrix array
   assign ecchmatrix[0][0] = 1;
   assign ecchmatrix[1][0] = 1;
   assign ecchmatrix[2][0] = 1;
   assign ecchmatrix[3][0] = 0;
   assign ecchmatrix[4][0] = 0;
   assign ecchmatrix[5][0] = 0;
   assign ecchmatrix[6][0] = 0;
   assign ecchmatrix[7][0] = 0;
   assign ecchmatrix[0][1] = 1;
   assign ecchmatrix[1][1] = 1;
   assign ecchmatrix[2][1] = 0;
   assign ecchmatrix[3][1] = 1;
   assign ecchmatrix[4][1] = 0;
   assign ecchmatrix[5][1] = 0;
   assign ecchmatrix[6][1] = 0;
   assign ecchmatrix[7][1] = 0;
   assign ecchmatrix[0][2] = 1;
   assign ecchmatrix[1][2] = 1;
   assign ecchmatrix[2][2] = 0;
   assign ecchmatrix[3][2] = 0;
   assign ecchmatrix[4][2] = 1;
   assign ecchmatrix[5][2] = 0;
   assign ecchmatrix[6][2] = 0;
   assign ecchmatrix[7][2] = 0;
   assign ecchmatrix[0][3] = 1;
   assign ecchmatrix[1][3] = 1;
   assign ecchmatrix[2][3] = 0;
   assign ecchmatrix[3][3] = 0;
   assign ecchmatrix[4][3] = 0;
   assign ecchmatrix[5][3] = 1;
   assign ecchmatrix[6][3] = 0;
   assign ecchmatrix[7][3] = 0;
   assign ecchmatrix[0][4] = 1;
   assign ecchmatrix[1][4] = 1;
   assign ecchmatrix[2][4] = 0;
   assign ecchmatrix[3][4] = 0;
   assign ecchmatrix[4][4] = 0;
   assign ecchmatrix[5][4] = 0;
   assign ecchmatrix[6][4] = 1;
   assign ecchmatrix[7][4] = 0;
   assign ecchmatrix[0][5] = 1;
   assign ecchmatrix[1][5] = 1;
   assign ecchmatrix[2][5] = 0;
   assign ecchmatrix[3][5] = 0;
   assign ecchmatrix[4][5] = 0;
   assign ecchmatrix[5][5] = 0;
   assign ecchmatrix[6][5] = 0;
   assign ecchmatrix[7][5] = 1;
   assign ecchmatrix[0][6] = 1;
   assign ecchmatrix[1][6] = 0;
   assign ecchmatrix[2][6] = 1;
   assign ecchmatrix[3][6] = 1;
   assign ecchmatrix[4][6] = 0;
   assign ecchmatrix[5][6] = 0;
   assign ecchmatrix[6][6] = 0;
   assign ecchmatrix[7][6] = 0;
   assign ecchmatrix[0][7] = 1;
   assign ecchmatrix[1][7] = 0;
   assign ecchmatrix[2][7] = 1;
   assign ecchmatrix[3][7] = 0;
   assign ecchmatrix[4][7] = 1;
   assign ecchmatrix[5][7] = 0;
   assign ecchmatrix[6][7] = 0;
   assign ecchmatrix[7][7] = 0;
   assign ecchmatrix[0][8] = 1;
   assign ecchmatrix[1][8] = 0;
   assign ecchmatrix[2][8] = 1;
   assign ecchmatrix[3][8] = 0;
   assign ecchmatrix[4][8] = 0;
   assign ecchmatrix[5][8] = 1;
   assign ecchmatrix[6][8] = 0;
   assign ecchmatrix[7][8] = 0;
   assign ecchmatrix[0][9] = 1;
   assign ecchmatrix[1][9] = 0;
   assign ecchmatrix[2][9] = 1;
   assign ecchmatrix[3][9] = 0;
   assign ecchmatrix[4][9] = 0;
   assign ecchmatrix[5][9] = 0;
   assign ecchmatrix[6][9] = 1;
   assign ecchmatrix[7][9] = 0;
   assign ecchmatrix[0][10] = 1;
   assign ecchmatrix[1][10] = 0;
   assign ecchmatrix[2][10] = 1;
   assign ecchmatrix[3][10] = 0;
   assign ecchmatrix[4][10] = 0;
   assign ecchmatrix[5][10] = 0;
   assign ecchmatrix[6][10] = 0;
   assign ecchmatrix[7][10] = 1;
   assign ecchmatrix[0][11] = 1;
   assign ecchmatrix[1][11] = 0;
   assign ecchmatrix[2][11] = 0;
   assign ecchmatrix[3][11] = 1;
   assign ecchmatrix[4][11] = 1;
   assign ecchmatrix[5][11] = 0;
   assign ecchmatrix[6][11] = 0;
   assign ecchmatrix[7][11] = 0;
   assign ecchmatrix[0][12] = 1;
   assign ecchmatrix[1][12] = 0;
   assign ecchmatrix[2][12] = 0;
   assign ecchmatrix[3][12] = 1;
   assign ecchmatrix[4][12] = 0;
   assign ecchmatrix[5][12] = 1;
   assign ecchmatrix[6][12] = 0;
   assign ecchmatrix[7][12] = 0;
   assign ecchmatrix[0][13] = 1;
   assign ecchmatrix[1][13] = 0;
   assign ecchmatrix[2][13] = 0;
   assign ecchmatrix[3][13] = 1;
   assign ecchmatrix[4][13] = 0;
   assign ecchmatrix[5][13] = 0;
   assign ecchmatrix[6][13] = 1;
   assign ecchmatrix[7][13] = 0;
   assign ecchmatrix[0][14] = 1;
   assign ecchmatrix[1][14] = 0;
   assign ecchmatrix[2][14] = 0;
   assign ecchmatrix[3][14] = 1;
   assign ecchmatrix[4][14] = 0;
   assign ecchmatrix[5][14] = 0;
   assign ecchmatrix[6][14] = 0;
   assign ecchmatrix[7][14] = 1;
   assign ecchmatrix[0][15] = 1;
   assign ecchmatrix[1][15] = 0;
   assign ecchmatrix[2][15] = 0;
   assign ecchmatrix[3][15] = 0;
   assign ecchmatrix[4][15] = 1;
   assign ecchmatrix[5][15] = 1;
   assign ecchmatrix[6][15] = 0;
   assign ecchmatrix[7][15] = 0;
   assign ecchmatrix[0][16] = 1;
   assign ecchmatrix[1][16] = 0;
   assign ecchmatrix[2][16] = 0;
   assign ecchmatrix[3][16] = 0;
   assign ecchmatrix[4][16] = 1;
   assign ecchmatrix[5][16] = 0;
   assign ecchmatrix[6][16] = 1;
   assign ecchmatrix[7][16] = 0;
   assign ecchmatrix[0][17] = 1;
   assign ecchmatrix[1][17] = 0;
   assign ecchmatrix[2][17] = 0;
   assign ecchmatrix[3][17] = 0;
   assign ecchmatrix[4][17] = 1;
   assign ecchmatrix[5][17] = 0;
   assign ecchmatrix[6][17] = 0;
   assign ecchmatrix[7][17] = 1;
   assign ecchmatrix[0][18] = 1;
   assign ecchmatrix[1][18] = 0;
   assign ecchmatrix[2][18] = 0;
   assign ecchmatrix[3][18] = 0;
   assign ecchmatrix[4][18] = 0;
   assign ecchmatrix[5][18] = 1;
   assign ecchmatrix[6][18] = 1;
   assign ecchmatrix[7][18] = 0;
   assign ecchmatrix[0][19] = 1;
   assign ecchmatrix[1][19] = 0;
   assign ecchmatrix[2][19] = 0;
   assign ecchmatrix[3][19] = 0;
   assign ecchmatrix[4][19] = 0;
   assign ecchmatrix[5][19] = 1;
   assign ecchmatrix[6][19] = 0;
   assign ecchmatrix[7][19] = 1;
   assign ecchmatrix[0][20] = 1;
   assign ecchmatrix[1][20] = 0;
   assign ecchmatrix[2][20] = 0;
   assign ecchmatrix[3][20] = 0;
   assign ecchmatrix[4][20] = 0;
   assign ecchmatrix[5][20] = 0;
   assign ecchmatrix[6][20] = 1;
   assign ecchmatrix[7][20] = 1;
   assign ecchmatrix[0][21] = 0;
   assign ecchmatrix[1][21] = 1;
   assign ecchmatrix[2][21] = 1;
   assign ecchmatrix[3][21] = 1;
   assign ecchmatrix[4][21] = 0;
   assign ecchmatrix[5][21] = 0;
   assign ecchmatrix[6][21] = 0;
   assign ecchmatrix[7][21] = 0;
   assign ecchmatrix[0][22] = 0;
   assign ecchmatrix[1][22] = 1;
   assign ecchmatrix[2][22] = 1;
   assign ecchmatrix[3][22] = 0;
   assign ecchmatrix[4][22] = 1;
   assign ecchmatrix[5][22] = 0;
   assign ecchmatrix[6][22] = 0;
   assign ecchmatrix[7][22] = 0;
   assign ecchmatrix[0][23] = 0;
   assign ecchmatrix[1][23] = 1;
   assign ecchmatrix[2][23] = 1;
   assign ecchmatrix[3][23] = 0;
   assign ecchmatrix[4][23] = 0;
   assign ecchmatrix[5][23] = 1;
   assign ecchmatrix[6][23] = 0;
   assign ecchmatrix[7][23] = 0;
   assign ecchmatrix[0][24] = 0;
   assign ecchmatrix[1][24] = 1;
   assign ecchmatrix[2][24] = 1;
   assign ecchmatrix[3][24] = 0;
   assign ecchmatrix[4][24] = 0;
   assign ecchmatrix[5][24] = 0;
   assign ecchmatrix[6][24] = 1;
   assign ecchmatrix[7][24] = 0;
   assign ecchmatrix[0][25] = 0;
   assign ecchmatrix[1][25] = 1;
   assign ecchmatrix[2][25] = 1;
   assign ecchmatrix[3][25] = 0;
   assign ecchmatrix[4][25] = 0;
   assign ecchmatrix[5][25] = 0;
   assign ecchmatrix[6][25] = 0;
   assign ecchmatrix[7][25] = 1;
   assign ecchmatrix[0][26] = 0;
   assign ecchmatrix[1][26] = 1;
   assign ecchmatrix[2][26] = 0;
   assign ecchmatrix[3][26] = 1;
   assign ecchmatrix[4][26] = 1;
   assign ecchmatrix[5][26] = 0;
   assign ecchmatrix[6][26] = 0;
   assign ecchmatrix[7][26] = 0;
   assign ecchmatrix[0][27] = 0;
   assign ecchmatrix[1][27] = 1;
   assign ecchmatrix[2][27] = 0;
   assign ecchmatrix[3][27] = 1;
   assign ecchmatrix[4][27] = 0;
   assign ecchmatrix[5][27] = 1;
   assign ecchmatrix[6][27] = 0;
   assign ecchmatrix[7][27] = 0;
   assign ecchmatrix[0][28] = 0;
   assign ecchmatrix[1][28] = 1;
   assign ecchmatrix[2][28] = 0;
   assign ecchmatrix[3][28] = 1;
   assign ecchmatrix[4][28] = 0;
   assign ecchmatrix[5][28] = 0;
   assign ecchmatrix[6][28] = 1;
   assign ecchmatrix[7][28] = 0;
   assign ecchmatrix[0][29] = 0;
   assign ecchmatrix[1][29] = 1;
   assign ecchmatrix[2][29] = 0;
   assign ecchmatrix[3][29] = 1;
   assign ecchmatrix[4][29] = 0;
   assign ecchmatrix[5][29] = 0;
   assign ecchmatrix[6][29] = 0;
   assign ecchmatrix[7][29] = 1;
   assign ecchmatrix[0][30] = 0;
   assign ecchmatrix[1][30] = 1;
   assign ecchmatrix[2][30] = 0;
   assign ecchmatrix[3][30] = 0;
   assign ecchmatrix[4][30] = 1;
   assign ecchmatrix[5][30] = 1;
   assign ecchmatrix[6][30] = 0;
   assign ecchmatrix[7][30] = 0;
   assign ecchmatrix[0][31] = 0;
   assign ecchmatrix[1][31] = 1;
   assign ecchmatrix[2][31] = 0;
   assign ecchmatrix[3][31] = 0;
   assign ecchmatrix[4][31] = 1;
   assign ecchmatrix[5][31] = 0;
   assign ecchmatrix[6][31] = 1;
   assign ecchmatrix[7][31] = 0;
   assign ecchmatrix[0][32] = 0;
   assign ecchmatrix[1][32] = 1;
   assign ecchmatrix[2][32] = 0;
   assign ecchmatrix[3][32] = 0;
   assign ecchmatrix[4][32] = 1;
   assign ecchmatrix[5][32] = 0;
   assign ecchmatrix[6][32] = 0;
   assign ecchmatrix[7][32] = 1;
   assign ecchmatrix[0][33] = 0;
   assign ecchmatrix[1][33] = 1;
   assign ecchmatrix[2][33] = 0;
   assign ecchmatrix[3][33] = 0;
   assign ecchmatrix[4][33] = 0;
   assign ecchmatrix[5][33] = 1;
   assign ecchmatrix[6][33] = 1;
   assign ecchmatrix[7][33] = 0;
   assign ecchmatrix[0][34] = 0;
   assign ecchmatrix[1][34] = 1;
   assign ecchmatrix[2][34] = 0;
   assign ecchmatrix[3][34] = 0;
   assign ecchmatrix[4][34] = 0;
   assign ecchmatrix[5][34] = 1;
   assign ecchmatrix[6][34] = 0;
   assign ecchmatrix[7][34] = 1;
   assign ecchmatrix[0][35] = 0;
   assign ecchmatrix[1][35] = 1;
   assign ecchmatrix[2][35] = 0;
   assign ecchmatrix[3][35] = 0;
   assign ecchmatrix[4][35] = 0;
   assign ecchmatrix[5][35] = 0;
   assign ecchmatrix[6][35] = 1;
   assign ecchmatrix[7][35] = 1;
   assign ecchmatrix[0][36] = 0;
   assign ecchmatrix[1][36] = 0;
   assign ecchmatrix[2][36] = 1;
   assign ecchmatrix[3][36] = 1;
   assign ecchmatrix[4][36] = 1;
   assign ecchmatrix[5][36] = 0;
   assign ecchmatrix[6][36] = 0;
   assign ecchmatrix[7][36] = 0;
   assign ecchmatrix[0][37] = 0;
   assign ecchmatrix[1][37] = 0;
   assign ecchmatrix[2][37] = 1;
   assign ecchmatrix[3][37] = 1;
   assign ecchmatrix[4][37] = 0;
   assign ecchmatrix[5][37] = 1;
   assign ecchmatrix[6][37] = 0;
   assign ecchmatrix[7][37] = 0;
   assign ecchmatrix[0][38] = 0;
   assign ecchmatrix[1][38] = 0;
   assign ecchmatrix[2][38] = 1;
   assign ecchmatrix[3][38] = 1;
   assign ecchmatrix[4][38] = 0;
   assign ecchmatrix[5][38] = 0;
   assign ecchmatrix[6][38] = 1;
   assign ecchmatrix[7][38] = 0;
   assign ecchmatrix[0][39] = 0;
   assign ecchmatrix[1][39] = 0;
   assign ecchmatrix[2][39] = 1;
   assign ecchmatrix[3][39] = 1;
   assign ecchmatrix[4][39] = 0;
   assign ecchmatrix[5][39] = 0;
   assign ecchmatrix[6][39] = 0;
   assign ecchmatrix[7][39] = 1;
   assign ecchmatrix[0][40] = 0;
   assign ecchmatrix[1][40] = 0;
   assign ecchmatrix[2][40] = 1;
   assign ecchmatrix[3][40] = 0;
   assign ecchmatrix[4][40] = 1;
   assign ecchmatrix[5][40] = 1;
   assign ecchmatrix[6][40] = 0;
   assign ecchmatrix[7][40] = 0;
   assign ecchmatrix[0][41] = 0;
   assign ecchmatrix[1][41] = 0;
   assign ecchmatrix[2][41] = 1;
   assign ecchmatrix[3][41] = 0;
   assign ecchmatrix[4][41] = 1;
   assign ecchmatrix[5][41] = 0;
   assign ecchmatrix[6][41] = 1;
   assign ecchmatrix[7][41] = 0;
   assign ecchmatrix[0][42] = 0;
   assign ecchmatrix[1][42] = 0;
   assign ecchmatrix[2][42] = 1;
   assign ecchmatrix[3][42] = 0;
   assign ecchmatrix[4][42] = 1;
   assign ecchmatrix[5][42] = 0;
   assign ecchmatrix[6][42] = 0;
   assign ecchmatrix[7][42] = 1;
   assign ecchmatrix[0][43] = 0;
   assign ecchmatrix[1][43] = 0;
   assign ecchmatrix[2][43] = 1;
   assign ecchmatrix[3][43] = 0;
   assign ecchmatrix[4][43] = 0;
   assign ecchmatrix[5][43] = 1;
   assign ecchmatrix[6][43] = 1;
   assign ecchmatrix[7][43] = 0;
   assign ecchmatrix[0][44] = 0;
   assign ecchmatrix[1][44] = 0;
   assign ecchmatrix[2][44] = 1;
   assign ecchmatrix[3][44] = 0;
   assign ecchmatrix[4][44] = 0;
   assign ecchmatrix[5][44] = 1;
   assign ecchmatrix[6][44] = 0;
   assign ecchmatrix[7][44] = 1;
   assign ecchmatrix[0][45] = 0;
   assign ecchmatrix[1][45] = 0;
   assign ecchmatrix[2][45] = 1;
   assign ecchmatrix[3][45] = 0;
   assign ecchmatrix[4][45] = 0;
   assign ecchmatrix[5][45] = 0;
   assign ecchmatrix[6][45] = 1;
   assign ecchmatrix[7][45] = 1;
   assign ecchmatrix[0][46] = 0;
   assign ecchmatrix[1][46] = 0;
   assign ecchmatrix[2][46] = 0;
   assign ecchmatrix[3][46] = 1;
   assign ecchmatrix[4][46] = 1;
   assign ecchmatrix[5][46] = 1;
   assign ecchmatrix[6][46] = 0;
   assign ecchmatrix[7][46] = 0;
   assign ecchmatrix[0][47] = 0;
   assign ecchmatrix[1][47] = 0;
   assign ecchmatrix[2][47] = 0;
   assign ecchmatrix[3][47] = 1;
   assign ecchmatrix[4][47] = 1;
   assign ecchmatrix[5][47] = 0;
   assign ecchmatrix[6][47] = 1;
   assign ecchmatrix[7][47] = 0;
   assign ecchmatrix[0][48] = 0;
   assign ecchmatrix[1][48] = 0;
   assign ecchmatrix[2][48] = 0;
   assign ecchmatrix[3][48] = 1;
   assign ecchmatrix[4][48] = 1;
   assign ecchmatrix[5][48] = 0;
   assign ecchmatrix[6][48] = 0;
   assign ecchmatrix[7][48] = 1;
   assign ecchmatrix[0][49] = 0;
   assign ecchmatrix[1][49] = 0;
   assign ecchmatrix[2][49] = 0;
   assign ecchmatrix[3][49] = 1;
   assign ecchmatrix[4][49] = 0;
   assign ecchmatrix[5][49] = 1;
   assign ecchmatrix[6][49] = 1;
   assign ecchmatrix[7][49] = 0;
   assign ecchmatrix[0][50] = 0;
   assign ecchmatrix[1][50] = 0;
   assign ecchmatrix[2][50] = 0;
   assign ecchmatrix[3][50] = 1;
   assign ecchmatrix[4][50] = 0;
   assign ecchmatrix[5][50] = 1;
   assign ecchmatrix[6][50] = 0;
   assign ecchmatrix[7][50] = 1;
   assign ecchmatrix[0][51] = 0;
   assign ecchmatrix[1][51] = 0;
   assign ecchmatrix[2][51] = 0;
   assign ecchmatrix[3][51] = 1;
   assign ecchmatrix[4][51] = 0;
   assign ecchmatrix[5][51] = 0;
   assign ecchmatrix[6][51] = 1;
   assign ecchmatrix[7][51] = 1;
   assign ecchmatrix[0][52] = 0;
   assign ecchmatrix[1][52] = 0;
   assign ecchmatrix[2][52] = 0;
   assign ecchmatrix[3][52] = 0;
   assign ecchmatrix[4][52] = 1;
   assign ecchmatrix[5][52] = 1;
   assign ecchmatrix[6][52] = 1;
   assign ecchmatrix[7][52] = 0;
   assign ecchmatrix[0][53] = 0;
   assign ecchmatrix[1][53] = 0;
   assign ecchmatrix[2][53] = 0;
   assign ecchmatrix[3][53] = 0;
   assign ecchmatrix[4][53] = 1;
   assign ecchmatrix[5][53] = 1;
   assign ecchmatrix[6][53] = 0;
   assign ecchmatrix[7][53] = 1;
   assign ecchmatrix[0][54] = 0;
   assign ecchmatrix[1][54] = 0;
   assign ecchmatrix[2][54] = 0;
   assign ecchmatrix[3][54] = 0;
   assign ecchmatrix[4][54] = 1;
   assign ecchmatrix[5][54] = 0;
   assign ecchmatrix[6][54] = 1;
   assign ecchmatrix[7][54] = 1;
   assign ecchmatrix[0][55] = 0;
   assign ecchmatrix[1][55] = 0;
   assign ecchmatrix[2][55] = 0;
   assign ecchmatrix[3][55] = 0;
   assign ecchmatrix[4][55] = 0;
   assign ecchmatrix[5][55] = 1;
   assign ecchmatrix[6][55] = 1;
   assign ecchmatrix[7][55] = 1;
   assign ecchmatrix[0][56] = 1;
   assign ecchmatrix[1][56] = 1;
   assign ecchmatrix[2][56] = 1;
   assign ecchmatrix[3][56] = 1;
   assign ecchmatrix[4][56] = 1;
   assign ecchmatrix[5][56] = 0;
   assign ecchmatrix[6][56] = 0;
   assign ecchmatrix[7][56] = 0;
   assign ecchmatrix[0][57] = 1;
   assign ecchmatrix[1][57] = 1;
   assign ecchmatrix[2][57] = 1;
   assign ecchmatrix[3][57] = 1;
   assign ecchmatrix[4][57] = 0;
   assign ecchmatrix[5][57] = 1;
   assign ecchmatrix[6][57] = 0;
   assign ecchmatrix[7][57] = 0;
   assign ecchmatrix[0][58] = 1;
   assign ecchmatrix[1][58] = 1;
   assign ecchmatrix[2][58] = 1;
   assign ecchmatrix[3][58] = 1;
   assign ecchmatrix[4][58] = 0;
   assign ecchmatrix[5][58] = 0;
   assign ecchmatrix[6][58] = 1;
   assign ecchmatrix[7][58] = 0;
   assign ecchmatrix[0][59] = 1;
   assign ecchmatrix[1][59] = 1;
   assign ecchmatrix[2][59] = 1;
   assign ecchmatrix[3][59] = 1;
   assign ecchmatrix[4][59] = 0;
   assign ecchmatrix[5][59] = 0;
   assign ecchmatrix[6][59] = 0;
   assign ecchmatrix[7][59] = 1;
   assign ecchmatrix[0][60] = 1;
   assign ecchmatrix[1][60] = 1;
   assign ecchmatrix[2][60] = 1;
   assign ecchmatrix[3][60] = 0;
   assign ecchmatrix[4][60] = 1;
   assign ecchmatrix[5][60] = 1;
   assign ecchmatrix[6][60] = 0;
   assign ecchmatrix[7][60] = 0;
   assign ecchmatrix[0][61] = 1;
   assign ecchmatrix[1][61] = 1;
   assign ecchmatrix[2][61] = 1;
   assign ecchmatrix[3][61] = 0;
   assign ecchmatrix[4][61] = 1;
   assign ecchmatrix[5][61] = 0;
   assign ecchmatrix[6][61] = 1;
   assign ecchmatrix[7][61] = 0;
   assign ecchmatrix[0][62] = 1;
   assign ecchmatrix[1][62] = 1;
   assign ecchmatrix[2][62] = 1;
   assign ecchmatrix[3][62] = 0;
   assign ecchmatrix[4][62] = 1;
   assign ecchmatrix[5][62] = 0;
   assign ecchmatrix[6][62] = 0;
   assign ecchmatrix[7][62] = 1;
   assign ecchmatrix[0][63] = 1;
   assign ecchmatrix[1][63] = 1;
   assign ecchmatrix[2][63] = 1;
   assign ecchmatrix[3][63] = 0;
   assign ecchmatrix[4][63] = 0;
   assign ecchmatrix[5][63] = 1;
   assign ecchmatrix[6][63] = 1;
   assign ecchmatrix[7][63] = 0;
   assign ecchmatrix[0][64] = 1;
   assign ecchmatrix[1][64] = 1;
   assign ecchmatrix[2][64] = 1;
   assign ecchmatrix[3][64] = 0;
   assign ecchmatrix[4][64] = 0;
   assign ecchmatrix[5][64] = 1;
   assign ecchmatrix[6][64] = 0;
   assign ecchmatrix[7][64] = 1;
   assign ecchmatrix[0][65] = 1;
   assign ecchmatrix[1][65] = 1;
   assign ecchmatrix[2][65] = 1;
   assign ecchmatrix[3][65] = 0;
   assign ecchmatrix[4][65] = 0;
   assign ecchmatrix[5][65] = 0;
   assign ecchmatrix[6][65] = 1;
   assign ecchmatrix[7][65] = 1;
   assign ecchmatrix[0][66] = 1;
   assign ecchmatrix[1][66] = 1;
   assign ecchmatrix[2][66] = 0;
   assign ecchmatrix[3][66] = 1;
   assign ecchmatrix[4][66] = 1;
   assign ecchmatrix[5][66] = 1;
   assign ecchmatrix[6][66] = 0;
   assign ecchmatrix[7][66] = 0;
   assign ecchmatrix[0][67] = 1;
   assign ecchmatrix[1][67] = 1;
   assign ecchmatrix[2][67] = 0;
   assign ecchmatrix[3][67] = 1;
   assign ecchmatrix[4][67] = 1;
   assign ecchmatrix[5][67] = 0;
   assign ecchmatrix[6][67] = 1;
   assign ecchmatrix[7][67] = 0;
   assign ecchmatrix[0][68] = 1;
   assign ecchmatrix[1][68] = 1;
   assign ecchmatrix[2][68] = 0;
   assign ecchmatrix[3][68] = 1;
   assign ecchmatrix[4][68] = 1;
   assign ecchmatrix[5][68] = 0;
   assign ecchmatrix[6][68] = 0;
   assign ecchmatrix[7][68] = 1;
   assign ecchmatrix[0][69] = 1;
   assign ecchmatrix[1][69] = 1;
   assign ecchmatrix[2][69] = 0;
   assign ecchmatrix[3][69] = 1;
   assign ecchmatrix[4][69] = 0;
   assign ecchmatrix[5][69] = 1;
   assign ecchmatrix[6][69] = 1;
   assign ecchmatrix[7][69] = 0;
   assign ecchmatrix[0][70] = 1;
   assign ecchmatrix[1][70] = 1;
   assign ecchmatrix[2][70] = 0;
   assign ecchmatrix[3][70] = 1;
   assign ecchmatrix[4][70] = 0;
   assign ecchmatrix[5][70] = 1;
   assign ecchmatrix[6][70] = 0;
   assign ecchmatrix[7][70] = 1;
   assign ecchmatrix[0][71] = 1;
   assign ecchmatrix[1][71] = 1;
   assign ecchmatrix[2][71] = 0;
   assign ecchmatrix[3][71] = 1;
   assign ecchmatrix[4][71] = 0;
   assign ecchmatrix[5][71] = 0;
   assign ecchmatrix[6][71] = 1;
   assign ecchmatrix[7][71] = 1;
   assign ecchmatrix[0][72] = 1;
   assign ecchmatrix[1][72] = 1;
   assign ecchmatrix[2][72] = 0;
   assign ecchmatrix[3][72] = 0;
   assign ecchmatrix[4][72] = 1;
   assign ecchmatrix[5][72] = 1;
   assign ecchmatrix[6][72] = 1;
   assign ecchmatrix[7][72] = 0;
   assign ecchmatrix[0][73] = 1;
   assign ecchmatrix[1][73] = 1;
   assign ecchmatrix[2][73] = 0;
   assign ecchmatrix[3][73] = 0;
   assign ecchmatrix[4][73] = 1;
   assign ecchmatrix[5][73] = 1;
   assign ecchmatrix[6][73] = 0;
   assign ecchmatrix[7][73] = 1;
   assign ecchmatrix[0][74] = 1;
   assign ecchmatrix[1][74] = 1;
   assign ecchmatrix[2][74] = 0;
   assign ecchmatrix[3][74] = 0;
   assign ecchmatrix[4][74] = 1;
   assign ecchmatrix[5][74] = 0;
   assign ecchmatrix[6][74] = 1;
   assign ecchmatrix[7][74] = 1;
   assign ecchmatrix[0][75] = 1;
   assign ecchmatrix[1][75] = 1;
   assign ecchmatrix[2][75] = 0;
   assign ecchmatrix[3][75] = 0;
   assign ecchmatrix[4][75] = 0;
   assign ecchmatrix[5][75] = 1;
   assign ecchmatrix[6][75] = 1;
   assign ecchmatrix[7][75] = 1;
   assign ecchmatrix[0][76] = 1;
   assign ecchmatrix[1][76] = 0;
   assign ecchmatrix[2][76] = 1;
   assign ecchmatrix[3][76] = 1;
   assign ecchmatrix[4][76] = 1;
   assign ecchmatrix[5][76] = 1;
   assign ecchmatrix[6][76] = 0;
   assign ecchmatrix[7][76] = 0;
   assign ecchmatrix[0][77] = 1;
   assign ecchmatrix[1][77] = 0;
   assign ecchmatrix[2][77] = 1;
   assign ecchmatrix[3][77] = 1;
   assign ecchmatrix[4][77] = 1;
   assign ecchmatrix[5][77] = 0;
   assign ecchmatrix[6][77] = 1;
   assign ecchmatrix[7][77] = 0;
   assign ecchmatrix[0][78] = 1;
   assign ecchmatrix[1][78] = 0;
   assign ecchmatrix[2][78] = 1;
   assign ecchmatrix[3][78] = 1;
   assign ecchmatrix[4][78] = 1;
   assign ecchmatrix[5][78] = 0;
   assign ecchmatrix[6][78] = 0;
   assign ecchmatrix[7][78] = 1;
   assign ecchmatrix[0][79] = 1;
   assign ecchmatrix[1][79] = 0;
   assign ecchmatrix[2][79] = 1;
   assign ecchmatrix[3][79] = 1;
   assign ecchmatrix[4][79] = 0;
   assign ecchmatrix[5][79] = 1;
   assign ecchmatrix[6][79] = 1;
   assign ecchmatrix[7][79] = 0;
   assign ecchmatrix[0][80] = 1;
   assign ecchmatrix[1][80] = 0;
   assign ecchmatrix[2][80] = 1;
   assign ecchmatrix[3][80] = 1;
   assign ecchmatrix[4][80] = 0;
   assign ecchmatrix[5][80] = 1;
   assign ecchmatrix[6][80] = 0;
   assign ecchmatrix[7][80] = 1;
   assign ecchmatrix[0][81] = 1;
   assign ecchmatrix[1][81] = 0;
   assign ecchmatrix[2][81] = 1;
   assign ecchmatrix[3][81] = 1;
   assign ecchmatrix[4][81] = 0;
   assign ecchmatrix[5][81] = 0;
   assign ecchmatrix[6][81] = 1;
   assign ecchmatrix[7][81] = 1;
   assign ecchmatrix[0][82] = 1;
   assign ecchmatrix[1][82] = 0;
   assign ecchmatrix[2][82] = 1;
   assign ecchmatrix[3][82] = 0;
   assign ecchmatrix[4][82] = 1;
   assign ecchmatrix[5][82] = 1;
   assign ecchmatrix[6][82] = 1;
   assign ecchmatrix[7][82] = 0;
   assign ecchmatrix[0][83] = 1;
   assign ecchmatrix[1][83] = 0;
   assign ecchmatrix[2][83] = 1;
   assign ecchmatrix[3][83] = 0;
   assign ecchmatrix[4][83] = 1;
   assign ecchmatrix[5][83] = 1;
   assign ecchmatrix[6][83] = 0;
   assign ecchmatrix[7][83] = 1;
   assign ecchmatrix[0][84] = 1;
   assign ecchmatrix[1][84] = 0;
   assign ecchmatrix[2][84] = 1;
   assign ecchmatrix[3][84] = 0;
   assign ecchmatrix[4][84] = 1;
   assign ecchmatrix[5][84] = 0;
   assign ecchmatrix[6][84] = 1;
   assign ecchmatrix[7][84] = 1;
   assign ecchmatrix[0][85] = 1;
   assign ecchmatrix[1][85] = 0;
   assign ecchmatrix[2][85] = 1;
   assign ecchmatrix[3][85] = 0;
   assign ecchmatrix[4][85] = 0;
   assign ecchmatrix[5][85] = 1;
   assign ecchmatrix[6][85] = 1;
   assign ecchmatrix[7][85] = 1;
   assign ecchmatrix[0][86] = 1;
   assign ecchmatrix[1][86] = 0;
   assign ecchmatrix[2][86] = 0;
   assign ecchmatrix[3][86] = 1;
   assign ecchmatrix[4][86] = 1;
   assign ecchmatrix[5][86] = 1;
   assign ecchmatrix[6][86] = 1;
   assign ecchmatrix[7][86] = 0;
   assign ecchmatrix[0][87] = 1;
   assign ecchmatrix[1][87] = 0;
   assign ecchmatrix[2][87] = 0;
   assign ecchmatrix[3][87] = 1;
   assign ecchmatrix[4][87] = 1;
   assign ecchmatrix[5][87] = 1;
   assign ecchmatrix[6][87] = 0;
   assign ecchmatrix[7][87] = 1;
   assign ecchmatrix[0][88] = 1;
   assign ecchmatrix[1][88] = 0;
   assign ecchmatrix[2][88] = 0;
   assign ecchmatrix[3][88] = 1;
   assign ecchmatrix[4][88] = 1;
   assign ecchmatrix[5][88] = 0;
   assign ecchmatrix[6][88] = 1;
   assign ecchmatrix[7][88] = 1;
   assign ecchmatrix[0][89] = 1;
   assign ecchmatrix[1][89] = 0;
   assign ecchmatrix[2][89] = 0;
   assign ecchmatrix[3][89] = 1;
   assign ecchmatrix[4][89] = 0;
   assign ecchmatrix[5][89] = 1;
   assign ecchmatrix[6][89] = 1;
   assign ecchmatrix[7][89] = 1;
   assign ecchmatrix[0][90] = 1;
   assign ecchmatrix[1][90] = 0;
   assign ecchmatrix[2][90] = 0;
   assign ecchmatrix[3][90] = 0;
   assign ecchmatrix[4][90] = 1;
   assign ecchmatrix[5][90] = 1;
   assign ecchmatrix[6][90] = 1;
   assign ecchmatrix[7][90] = 1;
   assign ecchmatrix[0][91] = 0;
   assign ecchmatrix[1][91] = 1;
   assign ecchmatrix[2][91] = 1;
   assign ecchmatrix[3][91] = 1;
   assign ecchmatrix[4][91] = 1;
   assign ecchmatrix[5][91] = 1;
   assign ecchmatrix[6][91] = 0;
   assign ecchmatrix[7][91] = 0;
   assign ecchmatrix[0][92] = 0;
   assign ecchmatrix[1][92] = 1;
   assign ecchmatrix[2][92] = 1;
   assign ecchmatrix[3][92] = 1;
   assign ecchmatrix[4][92] = 1;
   assign ecchmatrix[5][92] = 0;
   assign ecchmatrix[6][92] = 1;
   assign ecchmatrix[7][92] = 0;
   assign ecchmatrix[0][93] = 0;
   assign ecchmatrix[1][93] = 1;
   assign ecchmatrix[2][93] = 1;
   assign ecchmatrix[3][93] = 1;
   assign ecchmatrix[4][93] = 1;
   assign ecchmatrix[5][93] = 0;
   assign ecchmatrix[6][93] = 0;
   assign ecchmatrix[7][93] = 1;
   assign ecchmatrix[0][94] = 0;
   assign ecchmatrix[1][94] = 1;
   assign ecchmatrix[2][94] = 1;
   assign ecchmatrix[3][94] = 1;
   assign ecchmatrix[4][94] = 0;
   assign ecchmatrix[5][94] = 1;
   assign ecchmatrix[6][94] = 1;
   assign ecchmatrix[7][94] = 0;
   assign ecchmatrix[0][95] = 0;
   assign ecchmatrix[1][95] = 1;
   assign ecchmatrix[2][95] = 1;
   assign ecchmatrix[3][95] = 1;
   assign ecchmatrix[4][95] = 0;
   assign ecchmatrix[5][95] = 1;
   assign ecchmatrix[6][95] = 0;
   assign ecchmatrix[7][95] = 1;
   assign ecchmatrix[0][96] = 0;
   assign ecchmatrix[1][96] = 1;
   assign ecchmatrix[2][96] = 1;
   assign ecchmatrix[3][96] = 1;
   assign ecchmatrix[4][96] = 0;
   assign ecchmatrix[5][96] = 0;
   assign ecchmatrix[6][96] = 1;
   assign ecchmatrix[7][96] = 1;
   assign ecchmatrix[0][97] = 0;
   assign ecchmatrix[1][97] = 1;
   assign ecchmatrix[2][97] = 1;
   assign ecchmatrix[3][97] = 0;
   assign ecchmatrix[4][97] = 1;
   assign ecchmatrix[5][97] = 1;
   assign ecchmatrix[6][97] = 1;
   assign ecchmatrix[7][97] = 0;
   assign ecchmatrix[0][98] = 0;
   assign ecchmatrix[1][98] = 1;
   assign ecchmatrix[2][98] = 1;
   assign ecchmatrix[3][98] = 0;
   assign ecchmatrix[4][98] = 1;
   assign ecchmatrix[5][98] = 1;
   assign ecchmatrix[6][98] = 0;
   assign ecchmatrix[7][98] = 1;
   assign ecchmatrix[0][99] = 0;
   assign ecchmatrix[1][99] = 1;
   assign ecchmatrix[2][99] = 1;
   assign ecchmatrix[3][99] = 0;
   assign ecchmatrix[4][99] = 1;
   assign ecchmatrix[5][99] = 0;
   assign ecchmatrix[6][99] = 1;
   assign ecchmatrix[7][99] = 1;
   assign ecchmatrix[0][100] = 0;
   assign ecchmatrix[1][100] = 1;
   assign ecchmatrix[2][100] = 1;
   assign ecchmatrix[3][100] = 0;
   assign ecchmatrix[4][100] = 0;
   assign ecchmatrix[5][100] = 1;
   assign ecchmatrix[6][100] = 1;
   assign ecchmatrix[7][100] = 1;
   assign ecchmatrix[0][101] = 0;
   assign ecchmatrix[1][101] = 1;
   assign ecchmatrix[2][101] = 0;
   assign ecchmatrix[3][101] = 1;
   assign ecchmatrix[4][101] = 1;
   assign ecchmatrix[5][101] = 1;
   assign ecchmatrix[6][101] = 1;
   assign ecchmatrix[7][101] = 0;
   assign ecchmatrix[0][102] = 0;
   assign ecchmatrix[1][102] = 1;
   assign ecchmatrix[2][102] = 0;
   assign ecchmatrix[3][102] = 1;
   assign ecchmatrix[4][102] = 1;
   assign ecchmatrix[5][102] = 1;
   assign ecchmatrix[6][102] = 0;
   assign ecchmatrix[7][102] = 1;
   assign ecchmatrix[0][103] = 0;
   assign ecchmatrix[1][103] = 1;
   assign ecchmatrix[2][103] = 0;
   assign ecchmatrix[3][103] = 1;
   assign ecchmatrix[4][103] = 1;
   assign ecchmatrix[5][103] = 0;
   assign ecchmatrix[6][103] = 1;
   assign ecchmatrix[7][103] = 1;
   assign ecchmatrix[0][104] = 0;
   assign ecchmatrix[1][104] = 1;
   assign ecchmatrix[2][104] = 0;
   assign ecchmatrix[3][104] = 1;
   assign ecchmatrix[4][104] = 0;
   assign ecchmatrix[5][104] = 1;
   assign ecchmatrix[6][104] = 1;
   assign ecchmatrix[7][104] = 1;
   assign ecchmatrix[0][105] = 0;
   assign ecchmatrix[1][105] = 1;
   assign ecchmatrix[2][105] = 0;
   assign ecchmatrix[3][105] = 0;
   assign ecchmatrix[4][105] = 1;
   assign ecchmatrix[5][105] = 1;
   assign ecchmatrix[6][105] = 1;
   assign ecchmatrix[7][105] = 1;
   assign ecchmatrix[0][106] = 0;
   assign ecchmatrix[1][106] = 0;
   assign ecchmatrix[2][106] = 1;
   assign ecchmatrix[3][106] = 1;
   assign ecchmatrix[4][106] = 1;
   assign ecchmatrix[5][106] = 1;
   assign ecchmatrix[6][106] = 1;
   assign ecchmatrix[7][106] = 0;
   assign ecchmatrix[0][107] = 0;
   assign ecchmatrix[1][107] = 0;
   assign ecchmatrix[2][107] = 1;
   assign ecchmatrix[3][107] = 1;
   assign ecchmatrix[4][107] = 1;
   assign ecchmatrix[5][107] = 1;
   assign ecchmatrix[6][107] = 0;
   assign ecchmatrix[7][107] = 1;
   assign ecchmatrix[0][108] = 0;
   assign ecchmatrix[1][108] = 0;
   assign ecchmatrix[2][108] = 1;
   assign ecchmatrix[3][108] = 1;
   assign ecchmatrix[4][108] = 1;
   assign ecchmatrix[5][108] = 0;
   assign ecchmatrix[6][108] = 1;
   assign ecchmatrix[7][108] = 1;
   assign ecchmatrix[0][109] = 0;
   assign ecchmatrix[1][109] = 0;
   assign ecchmatrix[2][109] = 1;
   assign ecchmatrix[3][109] = 1;
   assign ecchmatrix[4][109] = 0;
   assign ecchmatrix[5][109] = 1;
   assign ecchmatrix[6][109] = 1;
   assign ecchmatrix[7][109] = 1;
   assign ecchmatrix[0][110] = 0;
   assign ecchmatrix[1][110] = 0;
   assign ecchmatrix[2][110] = 1;
   assign ecchmatrix[3][110] = 0;
   assign ecchmatrix[4][110] = 1;
   assign ecchmatrix[5][110] = 1;
   assign ecchmatrix[6][110] = 1;
   assign ecchmatrix[7][110] = 1;
   assign ecchmatrix[0][111] = 0;
   assign ecchmatrix[1][111] = 0;
   assign ecchmatrix[2][111] = 0;
   assign ecchmatrix[3][111] = 1;
   assign ecchmatrix[4][111] = 1;
   assign ecchmatrix[5][111] = 1;
   assign ecchmatrix[6][111] = 1;
   assign ecchmatrix[7][111] = 1;
   assign ecchmatrix[0][112] = 1;
   assign ecchmatrix[1][112] = 1;
   assign ecchmatrix[2][112] = 1;
   assign ecchmatrix[3][112] = 1;
   assign ecchmatrix[4][112] = 1;
   assign ecchmatrix[5][112] = 1;
   assign ecchmatrix[6][112] = 1;
   assign ecchmatrix[7][112] = 0;
   assign ecchmatrix[0][113] = 1;
   assign ecchmatrix[1][113] = 1;
   assign ecchmatrix[2][113] = 1;
   assign ecchmatrix[3][113] = 1;
   assign ecchmatrix[4][113] = 1;
   assign ecchmatrix[5][113] = 1;
   assign ecchmatrix[6][113] = 0;
   assign ecchmatrix[7][113] = 1;
   assign ecchmatrix[0][114] = 1;
   assign ecchmatrix[1][114] = 1;
   assign ecchmatrix[2][114] = 1;
   assign ecchmatrix[3][114] = 1;
   assign ecchmatrix[4][114] = 1;
   assign ecchmatrix[5][114] = 0;
   assign ecchmatrix[6][114] = 1;
   assign ecchmatrix[7][114] = 1;
   assign ecchmatrix[0][115] = 1;
   assign ecchmatrix[1][115] = 1;
   assign ecchmatrix[2][115] = 1;
   assign ecchmatrix[3][115] = 1;
   assign ecchmatrix[4][115] = 0;
   assign ecchmatrix[5][115] = 1;
   assign ecchmatrix[6][115] = 1;
   assign ecchmatrix[7][115] = 1;
   assign ecchmatrix[0][116] = 1;
   assign ecchmatrix[1][116] = 1;
   assign ecchmatrix[2][116] = 1;
   assign ecchmatrix[3][116] = 0;
   assign ecchmatrix[4][116] = 1;
   assign ecchmatrix[5][116] = 1;
   assign ecchmatrix[6][116] = 1;
   assign ecchmatrix[7][116] = 1;
   assign ecchmatrix[0][117] = 1;
   assign ecchmatrix[1][117] = 1;
   assign ecchmatrix[2][117] = 0;
   assign ecchmatrix[3][117] = 1;
   assign ecchmatrix[4][117] = 1;
   assign ecchmatrix[5][117] = 1;
   assign ecchmatrix[6][117] = 1;
   assign ecchmatrix[7][117] = 1;
   assign ecchmatrix[0][118] = 1;
   assign ecchmatrix[1][118] = 0;
   assign ecchmatrix[2][118] = 1;
   assign ecchmatrix[3][118] = 1;
   assign ecchmatrix[4][118] = 1;
   assign ecchmatrix[5][118] = 1;
   assign ecchmatrix[6][118] = 1;
   assign ecchmatrix[7][118] = 1;
   assign ecchmatrix[0][119] = 0;
   assign ecchmatrix[1][119] = 1;
   assign ecchmatrix[2][119] = 1;
   assign ecchmatrix[3][119] = 1;
   assign ecchmatrix[4][119] = 1;
   assign ecchmatrix[5][119] = 1;
   assign ecchmatrix[6][119] = 1;
   assign ecchmatrix[7][119] = 1;
endmodule

module ecc_calc_247 (din, eccout);

  localparam ECCDWIDTH = 247;
  localparam ECCWIDTH  = 9;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  wire [ECCDWIDTH-1:0]   ecchmatrix [0:ECCWIDTH-1];

 assign eccout[8] = ^(ecchmatrix[8]&din);
 assign eccout[7] = ^(ecchmatrix[7]&din);
 assign eccout[6] = ^(ecchmatrix[6]&din);
 assign eccout[5] = ^(ecchmatrix[5]&din);
 assign eccout[4] = ^(ecchmatrix[4]&din);
 assign eccout[3] = ^(ecchmatrix[3]&din);
 assign eccout[2] = ^(ecchmatrix[2]&din);
 assign eccout[1] = ^(ecchmatrix[1]&din);
 assign eccout[0] = ^(ecchmatrix[0]&din);
// assign ready = 1'b1;

// Generate the H Matrix in Perl

// Initialize the hmatrix array
   assign ecchmatrix[0][0] = 1;
   assign ecchmatrix[1][0] = 1;
   assign ecchmatrix[2][0] = 1;
   assign ecchmatrix[3][0] = 0;
   assign ecchmatrix[4][0] = 0;
   assign ecchmatrix[5][0] = 0;
   assign ecchmatrix[6][0] = 0;
   assign ecchmatrix[7][0] = 0;
   assign ecchmatrix[8][0] = 0;
   assign ecchmatrix[0][1] = 1;
   assign ecchmatrix[1][1] = 1;
   assign ecchmatrix[2][1] = 0;
   assign ecchmatrix[3][1] = 1;
   assign ecchmatrix[4][1] = 0;
   assign ecchmatrix[5][1] = 0;
   assign ecchmatrix[6][1] = 0;
   assign ecchmatrix[7][1] = 0;
   assign ecchmatrix[8][1] = 0;
   assign ecchmatrix[0][2] = 1;
   assign ecchmatrix[1][2] = 1;
   assign ecchmatrix[2][2] = 0;
   assign ecchmatrix[3][2] = 0;
   assign ecchmatrix[4][2] = 1;
   assign ecchmatrix[5][2] = 0;
   assign ecchmatrix[6][2] = 0;
   assign ecchmatrix[7][2] = 0;
   assign ecchmatrix[8][2] = 0;
   assign ecchmatrix[0][3] = 1;
   assign ecchmatrix[1][3] = 1;
   assign ecchmatrix[2][3] = 0;
   assign ecchmatrix[3][3] = 0;
   assign ecchmatrix[4][3] = 0;
   assign ecchmatrix[5][3] = 1;
   assign ecchmatrix[6][3] = 0;
   assign ecchmatrix[7][3] = 0;
   assign ecchmatrix[8][3] = 0;
   assign ecchmatrix[0][4] = 1;
   assign ecchmatrix[1][4] = 1;
   assign ecchmatrix[2][4] = 0;
   assign ecchmatrix[3][4] = 0;
   assign ecchmatrix[4][4] = 0;
   assign ecchmatrix[5][4] = 0;
   assign ecchmatrix[6][4] = 1;
   assign ecchmatrix[7][4] = 0;
   assign ecchmatrix[8][4] = 0;
   assign ecchmatrix[0][5] = 1;
   assign ecchmatrix[1][5] = 1;
   assign ecchmatrix[2][5] = 0;
   assign ecchmatrix[3][5] = 0;
   assign ecchmatrix[4][5] = 0;
   assign ecchmatrix[5][5] = 0;
   assign ecchmatrix[6][5] = 0;
   assign ecchmatrix[7][5] = 1;
   assign ecchmatrix[8][5] = 0;
   assign ecchmatrix[0][6] = 1;
   assign ecchmatrix[1][6] = 1;
   assign ecchmatrix[2][6] = 0;
   assign ecchmatrix[3][6] = 0;
   assign ecchmatrix[4][6] = 0;
   assign ecchmatrix[5][6] = 0;
   assign ecchmatrix[6][6] = 0;
   assign ecchmatrix[7][6] = 0;
   assign ecchmatrix[8][6] = 1;
   assign ecchmatrix[0][7] = 1;
   assign ecchmatrix[1][7] = 0;
   assign ecchmatrix[2][7] = 1;
   assign ecchmatrix[3][7] = 1;
   assign ecchmatrix[4][7] = 0;
   assign ecchmatrix[5][7] = 0;
   assign ecchmatrix[6][7] = 0;
   assign ecchmatrix[7][7] = 0;
   assign ecchmatrix[8][7] = 0;
   assign ecchmatrix[0][8] = 1;
   assign ecchmatrix[1][8] = 0;
   assign ecchmatrix[2][8] = 1;
   assign ecchmatrix[3][8] = 0;
   assign ecchmatrix[4][8] = 1;
   assign ecchmatrix[5][8] = 0;
   assign ecchmatrix[6][8] = 0;
   assign ecchmatrix[7][8] = 0;
   assign ecchmatrix[8][8] = 0;
   assign ecchmatrix[0][9] = 1;
   assign ecchmatrix[1][9] = 0;
   assign ecchmatrix[2][9] = 1;
   assign ecchmatrix[3][9] = 0;
   assign ecchmatrix[4][9] = 0;
   assign ecchmatrix[5][9] = 1;
   assign ecchmatrix[6][9] = 0;
   assign ecchmatrix[7][9] = 0;
   assign ecchmatrix[8][9] = 0;
   assign ecchmatrix[0][10] = 1;
   assign ecchmatrix[1][10] = 0;
   assign ecchmatrix[2][10] = 1;
   assign ecchmatrix[3][10] = 0;
   assign ecchmatrix[4][10] = 0;
   assign ecchmatrix[5][10] = 0;
   assign ecchmatrix[6][10] = 1;
   assign ecchmatrix[7][10] = 0;
   assign ecchmatrix[8][10] = 0;
   assign ecchmatrix[0][11] = 1;
   assign ecchmatrix[1][11] = 0;
   assign ecchmatrix[2][11] = 1;
   assign ecchmatrix[3][11] = 0;
   assign ecchmatrix[4][11] = 0;
   assign ecchmatrix[5][11] = 0;
   assign ecchmatrix[6][11] = 0;
   assign ecchmatrix[7][11] = 1;
   assign ecchmatrix[8][11] = 0;
   assign ecchmatrix[0][12] = 1;
   assign ecchmatrix[1][12] = 0;
   assign ecchmatrix[2][12] = 1;
   assign ecchmatrix[3][12] = 0;
   assign ecchmatrix[4][12] = 0;
   assign ecchmatrix[5][12] = 0;
   assign ecchmatrix[6][12] = 0;
   assign ecchmatrix[7][12] = 0;
   assign ecchmatrix[8][12] = 1;
   assign ecchmatrix[0][13] = 1;
   assign ecchmatrix[1][13] = 0;
   assign ecchmatrix[2][13] = 0;
   assign ecchmatrix[3][13] = 1;
   assign ecchmatrix[4][13] = 1;
   assign ecchmatrix[5][13] = 0;
   assign ecchmatrix[6][13] = 0;
   assign ecchmatrix[7][13] = 0;
   assign ecchmatrix[8][13] = 0;
   assign ecchmatrix[0][14] = 1;
   assign ecchmatrix[1][14] = 0;
   assign ecchmatrix[2][14] = 0;
   assign ecchmatrix[3][14] = 1;
   assign ecchmatrix[4][14] = 0;
   assign ecchmatrix[5][14] = 1;
   assign ecchmatrix[6][14] = 0;
   assign ecchmatrix[7][14] = 0;
   assign ecchmatrix[8][14] = 0;
   assign ecchmatrix[0][15] = 1;
   assign ecchmatrix[1][15] = 0;
   assign ecchmatrix[2][15] = 0;
   assign ecchmatrix[3][15] = 1;
   assign ecchmatrix[4][15] = 0;
   assign ecchmatrix[5][15] = 0;
   assign ecchmatrix[6][15] = 1;
   assign ecchmatrix[7][15] = 0;
   assign ecchmatrix[8][15] = 0;
   assign ecchmatrix[0][16] = 1;
   assign ecchmatrix[1][16] = 0;
   assign ecchmatrix[2][16] = 0;
   assign ecchmatrix[3][16] = 1;
   assign ecchmatrix[4][16] = 0;
   assign ecchmatrix[5][16] = 0;
   assign ecchmatrix[6][16] = 0;
   assign ecchmatrix[7][16] = 1;
   assign ecchmatrix[8][16] = 0;
   assign ecchmatrix[0][17] = 1;
   assign ecchmatrix[1][17] = 0;
   assign ecchmatrix[2][17] = 0;
   assign ecchmatrix[3][17] = 1;
   assign ecchmatrix[4][17] = 0;
   assign ecchmatrix[5][17] = 0;
   assign ecchmatrix[6][17] = 0;
   assign ecchmatrix[7][17] = 0;
   assign ecchmatrix[8][17] = 1;
   assign ecchmatrix[0][18] = 1;
   assign ecchmatrix[1][18] = 0;
   assign ecchmatrix[2][18] = 0;
   assign ecchmatrix[3][18] = 0;
   assign ecchmatrix[4][18] = 1;
   assign ecchmatrix[5][18] = 1;
   assign ecchmatrix[6][18] = 0;
   assign ecchmatrix[7][18] = 0;
   assign ecchmatrix[8][18] = 0;
   assign ecchmatrix[0][19] = 1;
   assign ecchmatrix[1][19] = 0;
   assign ecchmatrix[2][19] = 0;
   assign ecchmatrix[3][19] = 0;
   assign ecchmatrix[4][19] = 1;
   assign ecchmatrix[5][19] = 0;
   assign ecchmatrix[6][19] = 1;
   assign ecchmatrix[7][19] = 0;
   assign ecchmatrix[8][19] = 0;
   assign ecchmatrix[0][20] = 1;
   assign ecchmatrix[1][20] = 0;
   assign ecchmatrix[2][20] = 0;
   assign ecchmatrix[3][20] = 0;
   assign ecchmatrix[4][20] = 1;
   assign ecchmatrix[5][20] = 0;
   assign ecchmatrix[6][20] = 0;
   assign ecchmatrix[7][20] = 1;
   assign ecchmatrix[8][20] = 0;
   assign ecchmatrix[0][21] = 1;
   assign ecchmatrix[1][21] = 0;
   assign ecchmatrix[2][21] = 0;
   assign ecchmatrix[3][21] = 0;
   assign ecchmatrix[4][21] = 1;
   assign ecchmatrix[5][21] = 0;
   assign ecchmatrix[6][21] = 0;
   assign ecchmatrix[7][21] = 0;
   assign ecchmatrix[8][21] = 1;
   assign ecchmatrix[0][22] = 1;
   assign ecchmatrix[1][22] = 0;
   assign ecchmatrix[2][22] = 0;
   assign ecchmatrix[3][22] = 0;
   assign ecchmatrix[4][22] = 0;
   assign ecchmatrix[5][22] = 1;
   assign ecchmatrix[6][22] = 1;
   assign ecchmatrix[7][22] = 0;
   assign ecchmatrix[8][22] = 0;
   assign ecchmatrix[0][23] = 1;
   assign ecchmatrix[1][23] = 0;
   assign ecchmatrix[2][23] = 0;
   assign ecchmatrix[3][23] = 0;
   assign ecchmatrix[4][23] = 0;
   assign ecchmatrix[5][23] = 1;
   assign ecchmatrix[6][23] = 0;
   assign ecchmatrix[7][23] = 1;
   assign ecchmatrix[8][23] = 0;
   assign ecchmatrix[0][24] = 1;
   assign ecchmatrix[1][24] = 0;
   assign ecchmatrix[2][24] = 0;
   assign ecchmatrix[3][24] = 0;
   assign ecchmatrix[4][24] = 0;
   assign ecchmatrix[5][24] = 1;
   assign ecchmatrix[6][24] = 0;
   assign ecchmatrix[7][24] = 0;
   assign ecchmatrix[8][24] = 1;
   assign ecchmatrix[0][25] = 1;
   assign ecchmatrix[1][25] = 0;
   assign ecchmatrix[2][25] = 0;
   assign ecchmatrix[3][25] = 0;
   assign ecchmatrix[4][25] = 0;
   assign ecchmatrix[5][25] = 0;
   assign ecchmatrix[6][25] = 1;
   assign ecchmatrix[7][25] = 1;
   assign ecchmatrix[8][25] = 0;
   assign ecchmatrix[0][26] = 1;
   assign ecchmatrix[1][26] = 0;
   assign ecchmatrix[2][26] = 0;
   assign ecchmatrix[3][26] = 0;
   assign ecchmatrix[4][26] = 0;
   assign ecchmatrix[5][26] = 0;
   assign ecchmatrix[6][26] = 1;
   assign ecchmatrix[7][26] = 0;
   assign ecchmatrix[8][26] = 1;
   assign ecchmatrix[0][27] = 1;
   assign ecchmatrix[1][27] = 0;
   assign ecchmatrix[2][27] = 0;
   assign ecchmatrix[3][27] = 0;
   assign ecchmatrix[4][27] = 0;
   assign ecchmatrix[5][27] = 0;
   assign ecchmatrix[6][27] = 0;
   assign ecchmatrix[7][27] = 1;
   assign ecchmatrix[8][27] = 1;
   assign ecchmatrix[0][28] = 0;
   assign ecchmatrix[1][28] = 1;
   assign ecchmatrix[2][28] = 1;
   assign ecchmatrix[3][28] = 1;
   assign ecchmatrix[4][28] = 0;
   assign ecchmatrix[5][28] = 0;
   assign ecchmatrix[6][28] = 0;
   assign ecchmatrix[7][28] = 0;
   assign ecchmatrix[8][28] = 0;
   assign ecchmatrix[0][29] = 0;
   assign ecchmatrix[1][29] = 1;
   assign ecchmatrix[2][29] = 1;
   assign ecchmatrix[3][29] = 0;
   assign ecchmatrix[4][29] = 1;
   assign ecchmatrix[5][29] = 0;
   assign ecchmatrix[6][29] = 0;
   assign ecchmatrix[7][29] = 0;
   assign ecchmatrix[8][29] = 0;
   assign ecchmatrix[0][30] = 0;
   assign ecchmatrix[1][30] = 1;
   assign ecchmatrix[2][30] = 1;
   assign ecchmatrix[3][30] = 0;
   assign ecchmatrix[4][30] = 0;
   assign ecchmatrix[5][30] = 1;
   assign ecchmatrix[6][30] = 0;
   assign ecchmatrix[7][30] = 0;
   assign ecchmatrix[8][30] = 0;
   assign ecchmatrix[0][31] = 0;
   assign ecchmatrix[1][31] = 1;
   assign ecchmatrix[2][31] = 1;
   assign ecchmatrix[3][31] = 0;
   assign ecchmatrix[4][31] = 0;
   assign ecchmatrix[5][31] = 0;
   assign ecchmatrix[6][31] = 1;
   assign ecchmatrix[7][31] = 0;
   assign ecchmatrix[8][31] = 0;
   assign ecchmatrix[0][32] = 0;
   assign ecchmatrix[1][32] = 1;
   assign ecchmatrix[2][32] = 1;
   assign ecchmatrix[3][32] = 0;
   assign ecchmatrix[4][32] = 0;
   assign ecchmatrix[5][32] = 0;
   assign ecchmatrix[6][32] = 0;
   assign ecchmatrix[7][32] = 1;
   assign ecchmatrix[8][32] = 0;
   assign ecchmatrix[0][33] = 0;
   assign ecchmatrix[1][33] = 1;
   assign ecchmatrix[2][33] = 1;
   assign ecchmatrix[3][33] = 0;
   assign ecchmatrix[4][33] = 0;
   assign ecchmatrix[5][33] = 0;
   assign ecchmatrix[6][33] = 0;
   assign ecchmatrix[7][33] = 0;
   assign ecchmatrix[8][33] = 1;
   assign ecchmatrix[0][34] = 0;
   assign ecchmatrix[1][34] = 1;
   assign ecchmatrix[2][34] = 0;
   assign ecchmatrix[3][34] = 1;
   assign ecchmatrix[4][34] = 1;
   assign ecchmatrix[5][34] = 0;
   assign ecchmatrix[6][34] = 0;
   assign ecchmatrix[7][34] = 0;
   assign ecchmatrix[8][34] = 0;
   assign ecchmatrix[0][35] = 0;
   assign ecchmatrix[1][35] = 1;
   assign ecchmatrix[2][35] = 0;
   assign ecchmatrix[3][35] = 1;
   assign ecchmatrix[4][35] = 0;
   assign ecchmatrix[5][35] = 1;
   assign ecchmatrix[6][35] = 0;
   assign ecchmatrix[7][35] = 0;
   assign ecchmatrix[8][35] = 0;
   assign ecchmatrix[0][36] = 0;
   assign ecchmatrix[1][36] = 1;
   assign ecchmatrix[2][36] = 0;
   assign ecchmatrix[3][36] = 1;
   assign ecchmatrix[4][36] = 0;
   assign ecchmatrix[5][36] = 0;
   assign ecchmatrix[6][36] = 1;
   assign ecchmatrix[7][36] = 0;
   assign ecchmatrix[8][36] = 0;
   assign ecchmatrix[0][37] = 0;
   assign ecchmatrix[1][37] = 1;
   assign ecchmatrix[2][37] = 0;
   assign ecchmatrix[3][37] = 1;
   assign ecchmatrix[4][37] = 0;
   assign ecchmatrix[5][37] = 0;
   assign ecchmatrix[6][37] = 0;
   assign ecchmatrix[7][37] = 1;
   assign ecchmatrix[8][37] = 0;
   assign ecchmatrix[0][38] = 0;
   assign ecchmatrix[1][38] = 1;
   assign ecchmatrix[2][38] = 0;
   assign ecchmatrix[3][38] = 1;
   assign ecchmatrix[4][38] = 0;
   assign ecchmatrix[5][38] = 0;
   assign ecchmatrix[6][38] = 0;
   assign ecchmatrix[7][38] = 0;
   assign ecchmatrix[8][38] = 1;
   assign ecchmatrix[0][39] = 0;
   assign ecchmatrix[1][39] = 1;
   assign ecchmatrix[2][39] = 0;
   assign ecchmatrix[3][39] = 0;
   assign ecchmatrix[4][39] = 1;
   assign ecchmatrix[5][39] = 1;
   assign ecchmatrix[6][39] = 0;
   assign ecchmatrix[7][39] = 0;
   assign ecchmatrix[8][39] = 0;
   assign ecchmatrix[0][40] = 0;
   assign ecchmatrix[1][40] = 1;
   assign ecchmatrix[2][40] = 0;
   assign ecchmatrix[3][40] = 0;
   assign ecchmatrix[4][40] = 1;
   assign ecchmatrix[5][40] = 0;
   assign ecchmatrix[6][40] = 1;
   assign ecchmatrix[7][40] = 0;
   assign ecchmatrix[8][40] = 0;
   assign ecchmatrix[0][41] = 0;
   assign ecchmatrix[1][41] = 1;
   assign ecchmatrix[2][41] = 0;
   assign ecchmatrix[3][41] = 0;
   assign ecchmatrix[4][41] = 1;
   assign ecchmatrix[5][41] = 0;
   assign ecchmatrix[6][41] = 0;
   assign ecchmatrix[7][41] = 1;
   assign ecchmatrix[8][41] = 0;
   assign ecchmatrix[0][42] = 0;
   assign ecchmatrix[1][42] = 1;
   assign ecchmatrix[2][42] = 0;
   assign ecchmatrix[3][42] = 0;
   assign ecchmatrix[4][42] = 1;
   assign ecchmatrix[5][42] = 0;
   assign ecchmatrix[6][42] = 0;
   assign ecchmatrix[7][42] = 0;
   assign ecchmatrix[8][42] = 1;
   assign ecchmatrix[0][43] = 0;
   assign ecchmatrix[1][43] = 1;
   assign ecchmatrix[2][43] = 0;
   assign ecchmatrix[3][43] = 0;
   assign ecchmatrix[4][43] = 0;
   assign ecchmatrix[5][43] = 1;
   assign ecchmatrix[6][43] = 1;
   assign ecchmatrix[7][43] = 0;
   assign ecchmatrix[8][43] = 0;
   assign ecchmatrix[0][44] = 0;
   assign ecchmatrix[1][44] = 1;
   assign ecchmatrix[2][44] = 0;
   assign ecchmatrix[3][44] = 0;
   assign ecchmatrix[4][44] = 0;
   assign ecchmatrix[5][44] = 1;
   assign ecchmatrix[6][44] = 0;
   assign ecchmatrix[7][44] = 1;
   assign ecchmatrix[8][44] = 0;
   assign ecchmatrix[0][45] = 0;
   assign ecchmatrix[1][45] = 1;
   assign ecchmatrix[2][45] = 0;
   assign ecchmatrix[3][45] = 0;
   assign ecchmatrix[4][45] = 0;
   assign ecchmatrix[5][45] = 1;
   assign ecchmatrix[6][45] = 0;
   assign ecchmatrix[7][45] = 0;
   assign ecchmatrix[8][45] = 1;
   assign ecchmatrix[0][46] = 0;
   assign ecchmatrix[1][46] = 1;
   assign ecchmatrix[2][46] = 0;
   assign ecchmatrix[3][46] = 0;
   assign ecchmatrix[4][46] = 0;
   assign ecchmatrix[5][46] = 0;
   assign ecchmatrix[6][46] = 1;
   assign ecchmatrix[7][46] = 1;
   assign ecchmatrix[8][46] = 0;
   assign ecchmatrix[0][47] = 0;
   assign ecchmatrix[1][47] = 1;
   assign ecchmatrix[2][47] = 0;
   assign ecchmatrix[3][47] = 0;
   assign ecchmatrix[4][47] = 0;
   assign ecchmatrix[5][47] = 0;
   assign ecchmatrix[6][47] = 1;
   assign ecchmatrix[7][47] = 0;
   assign ecchmatrix[8][47] = 1;
   assign ecchmatrix[0][48] = 0;
   assign ecchmatrix[1][48] = 1;
   assign ecchmatrix[2][48] = 0;
   assign ecchmatrix[3][48] = 0;
   assign ecchmatrix[4][48] = 0;
   assign ecchmatrix[5][48] = 0;
   assign ecchmatrix[6][48] = 0;
   assign ecchmatrix[7][48] = 1;
   assign ecchmatrix[8][48] = 1;
   assign ecchmatrix[0][49] = 0;
   assign ecchmatrix[1][49] = 0;
   assign ecchmatrix[2][49] = 1;
   assign ecchmatrix[3][49] = 1;
   assign ecchmatrix[4][49] = 1;
   assign ecchmatrix[5][49] = 0;
   assign ecchmatrix[6][49] = 0;
   assign ecchmatrix[7][49] = 0;
   assign ecchmatrix[8][49] = 0;
   assign ecchmatrix[0][50] = 0;
   assign ecchmatrix[1][50] = 0;
   assign ecchmatrix[2][50] = 1;
   assign ecchmatrix[3][50] = 1;
   assign ecchmatrix[4][50] = 0;
   assign ecchmatrix[5][50] = 1;
   assign ecchmatrix[6][50] = 0;
   assign ecchmatrix[7][50] = 0;
   assign ecchmatrix[8][50] = 0;
   assign ecchmatrix[0][51] = 0;
   assign ecchmatrix[1][51] = 0;
   assign ecchmatrix[2][51] = 1;
   assign ecchmatrix[3][51] = 1;
   assign ecchmatrix[4][51] = 0;
   assign ecchmatrix[5][51] = 0;
   assign ecchmatrix[6][51] = 1;
   assign ecchmatrix[7][51] = 0;
   assign ecchmatrix[8][51] = 0;
   assign ecchmatrix[0][52] = 0;
   assign ecchmatrix[1][52] = 0;
   assign ecchmatrix[2][52] = 1;
   assign ecchmatrix[3][52] = 1;
   assign ecchmatrix[4][52] = 0;
   assign ecchmatrix[5][52] = 0;
   assign ecchmatrix[6][52] = 0;
   assign ecchmatrix[7][52] = 1;
   assign ecchmatrix[8][52] = 0;
   assign ecchmatrix[0][53] = 0;
   assign ecchmatrix[1][53] = 0;
   assign ecchmatrix[2][53] = 1;
   assign ecchmatrix[3][53] = 1;
   assign ecchmatrix[4][53] = 0;
   assign ecchmatrix[5][53] = 0;
   assign ecchmatrix[6][53] = 0;
   assign ecchmatrix[7][53] = 0;
   assign ecchmatrix[8][53] = 1;
   assign ecchmatrix[0][54] = 0;
   assign ecchmatrix[1][54] = 0;
   assign ecchmatrix[2][54] = 1;
   assign ecchmatrix[3][54] = 0;
   assign ecchmatrix[4][54] = 1;
   assign ecchmatrix[5][54] = 1;
   assign ecchmatrix[6][54] = 0;
   assign ecchmatrix[7][54] = 0;
   assign ecchmatrix[8][54] = 0;
   assign ecchmatrix[0][55] = 0;
   assign ecchmatrix[1][55] = 0;
   assign ecchmatrix[2][55] = 1;
   assign ecchmatrix[3][55] = 0;
   assign ecchmatrix[4][55] = 1;
   assign ecchmatrix[5][55] = 0;
   assign ecchmatrix[6][55] = 1;
   assign ecchmatrix[7][55] = 0;
   assign ecchmatrix[8][55] = 0;
   assign ecchmatrix[0][56] = 0;
   assign ecchmatrix[1][56] = 0;
   assign ecchmatrix[2][56] = 1;
   assign ecchmatrix[3][56] = 0;
   assign ecchmatrix[4][56] = 1;
   assign ecchmatrix[5][56] = 0;
   assign ecchmatrix[6][56] = 0;
   assign ecchmatrix[7][56] = 1;
   assign ecchmatrix[8][56] = 0;
   assign ecchmatrix[0][57] = 0;
   assign ecchmatrix[1][57] = 0;
   assign ecchmatrix[2][57] = 1;
   assign ecchmatrix[3][57] = 0;
   assign ecchmatrix[4][57] = 1;
   assign ecchmatrix[5][57] = 0;
   assign ecchmatrix[6][57] = 0;
   assign ecchmatrix[7][57] = 0;
   assign ecchmatrix[8][57] = 1;
   assign ecchmatrix[0][58] = 0;
   assign ecchmatrix[1][58] = 0;
   assign ecchmatrix[2][58] = 1;
   assign ecchmatrix[3][58] = 0;
   assign ecchmatrix[4][58] = 0;
   assign ecchmatrix[5][58] = 1;
   assign ecchmatrix[6][58] = 1;
   assign ecchmatrix[7][58] = 0;
   assign ecchmatrix[8][58] = 0;
   assign ecchmatrix[0][59] = 0;
   assign ecchmatrix[1][59] = 0;
   assign ecchmatrix[2][59] = 1;
   assign ecchmatrix[3][59] = 0;
   assign ecchmatrix[4][59] = 0;
   assign ecchmatrix[5][59] = 1;
   assign ecchmatrix[6][59] = 0;
   assign ecchmatrix[7][59] = 1;
   assign ecchmatrix[8][59] = 0;
   assign ecchmatrix[0][60] = 0;
   assign ecchmatrix[1][60] = 0;
   assign ecchmatrix[2][60] = 1;
   assign ecchmatrix[3][60] = 0;
   assign ecchmatrix[4][60] = 0;
   assign ecchmatrix[5][60] = 1;
   assign ecchmatrix[6][60] = 0;
   assign ecchmatrix[7][60] = 0;
   assign ecchmatrix[8][60] = 1;
   assign ecchmatrix[0][61] = 0;
   assign ecchmatrix[1][61] = 0;
   assign ecchmatrix[2][61] = 1;
   assign ecchmatrix[3][61] = 0;
   assign ecchmatrix[4][61] = 0;
   assign ecchmatrix[5][61] = 0;
   assign ecchmatrix[6][61] = 1;
   assign ecchmatrix[7][61] = 1;
   assign ecchmatrix[8][61] = 0;
   assign ecchmatrix[0][62] = 0;
   assign ecchmatrix[1][62] = 0;
   assign ecchmatrix[2][62] = 1;
   assign ecchmatrix[3][62] = 0;
   assign ecchmatrix[4][62] = 0;
   assign ecchmatrix[5][62] = 0;
   assign ecchmatrix[6][62] = 1;
   assign ecchmatrix[7][62] = 0;
   assign ecchmatrix[8][62] = 1;
   assign ecchmatrix[0][63] = 0;
   assign ecchmatrix[1][63] = 0;
   assign ecchmatrix[2][63] = 1;
   assign ecchmatrix[3][63] = 0;
   assign ecchmatrix[4][63] = 0;
   assign ecchmatrix[5][63] = 0;
   assign ecchmatrix[6][63] = 0;
   assign ecchmatrix[7][63] = 1;
   assign ecchmatrix[8][63] = 1;
   assign ecchmatrix[0][64] = 0;
   assign ecchmatrix[1][64] = 0;
   assign ecchmatrix[2][64] = 0;
   assign ecchmatrix[3][64] = 1;
   assign ecchmatrix[4][64] = 1;
   assign ecchmatrix[5][64] = 1;
   assign ecchmatrix[6][64] = 0;
   assign ecchmatrix[7][64] = 0;
   assign ecchmatrix[8][64] = 0;
   assign ecchmatrix[0][65] = 0;
   assign ecchmatrix[1][65] = 0;
   assign ecchmatrix[2][65] = 0;
   assign ecchmatrix[3][65] = 1;
   assign ecchmatrix[4][65] = 1;
   assign ecchmatrix[5][65] = 0;
   assign ecchmatrix[6][65] = 1;
   assign ecchmatrix[7][65] = 0;
   assign ecchmatrix[8][65] = 0;
   assign ecchmatrix[0][66] = 0;
   assign ecchmatrix[1][66] = 0;
   assign ecchmatrix[2][66] = 0;
   assign ecchmatrix[3][66] = 1;
   assign ecchmatrix[4][66] = 1;
   assign ecchmatrix[5][66] = 0;
   assign ecchmatrix[6][66] = 0;
   assign ecchmatrix[7][66] = 1;
   assign ecchmatrix[8][66] = 0;
   assign ecchmatrix[0][67] = 0;
   assign ecchmatrix[1][67] = 0;
   assign ecchmatrix[2][67] = 0;
   assign ecchmatrix[3][67] = 1;
   assign ecchmatrix[4][67] = 1;
   assign ecchmatrix[5][67] = 0;
   assign ecchmatrix[6][67] = 0;
   assign ecchmatrix[7][67] = 0;
   assign ecchmatrix[8][67] = 1;
   assign ecchmatrix[0][68] = 0;
   assign ecchmatrix[1][68] = 0;
   assign ecchmatrix[2][68] = 0;
   assign ecchmatrix[3][68] = 1;
   assign ecchmatrix[4][68] = 0;
   assign ecchmatrix[5][68] = 1;
   assign ecchmatrix[6][68] = 1;
   assign ecchmatrix[7][68] = 0;
   assign ecchmatrix[8][68] = 0;
   assign ecchmatrix[0][69] = 0;
   assign ecchmatrix[1][69] = 0;
   assign ecchmatrix[2][69] = 0;
   assign ecchmatrix[3][69] = 1;
   assign ecchmatrix[4][69] = 0;
   assign ecchmatrix[5][69] = 1;
   assign ecchmatrix[6][69] = 0;
   assign ecchmatrix[7][69] = 1;
   assign ecchmatrix[8][69] = 0;
   assign ecchmatrix[0][70] = 0;
   assign ecchmatrix[1][70] = 0;
   assign ecchmatrix[2][70] = 0;
   assign ecchmatrix[3][70] = 1;
   assign ecchmatrix[4][70] = 0;
   assign ecchmatrix[5][70] = 1;
   assign ecchmatrix[6][70] = 0;
   assign ecchmatrix[7][70] = 0;
   assign ecchmatrix[8][70] = 1;
   assign ecchmatrix[0][71] = 0;
   assign ecchmatrix[1][71] = 0;
   assign ecchmatrix[2][71] = 0;
   assign ecchmatrix[3][71] = 1;
   assign ecchmatrix[4][71] = 0;
   assign ecchmatrix[5][71] = 0;
   assign ecchmatrix[6][71] = 1;
   assign ecchmatrix[7][71] = 1;
   assign ecchmatrix[8][71] = 0;
   assign ecchmatrix[0][72] = 0;
   assign ecchmatrix[1][72] = 0;
   assign ecchmatrix[2][72] = 0;
   assign ecchmatrix[3][72] = 1;
   assign ecchmatrix[4][72] = 0;
   assign ecchmatrix[5][72] = 0;
   assign ecchmatrix[6][72] = 1;
   assign ecchmatrix[7][72] = 0;
   assign ecchmatrix[8][72] = 1;
   assign ecchmatrix[0][73] = 0;
   assign ecchmatrix[1][73] = 0;
   assign ecchmatrix[2][73] = 0;
   assign ecchmatrix[3][73] = 1;
   assign ecchmatrix[4][73] = 0;
   assign ecchmatrix[5][73] = 0;
   assign ecchmatrix[6][73] = 0;
   assign ecchmatrix[7][73] = 1;
   assign ecchmatrix[8][73] = 1;
   assign ecchmatrix[0][74] = 0;
   assign ecchmatrix[1][74] = 0;
   assign ecchmatrix[2][74] = 0;
   assign ecchmatrix[3][74] = 0;
   assign ecchmatrix[4][74] = 1;
   assign ecchmatrix[5][74] = 1;
   assign ecchmatrix[6][74] = 1;
   assign ecchmatrix[7][74] = 0;
   assign ecchmatrix[8][74] = 0;
   assign ecchmatrix[0][75] = 0;
   assign ecchmatrix[1][75] = 0;
   assign ecchmatrix[2][75] = 0;
   assign ecchmatrix[3][75] = 0;
   assign ecchmatrix[4][75] = 1;
   assign ecchmatrix[5][75] = 1;
   assign ecchmatrix[6][75] = 0;
   assign ecchmatrix[7][75] = 1;
   assign ecchmatrix[8][75] = 0;
   assign ecchmatrix[0][76] = 0;
   assign ecchmatrix[1][76] = 0;
   assign ecchmatrix[2][76] = 0;
   assign ecchmatrix[3][76] = 0;
   assign ecchmatrix[4][76] = 1;
   assign ecchmatrix[5][76] = 1;
   assign ecchmatrix[6][76] = 0;
   assign ecchmatrix[7][76] = 0;
   assign ecchmatrix[8][76] = 1;
   assign ecchmatrix[0][77] = 0;
   assign ecchmatrix[1][77] = 0;
   assign ecchmatrix[2][77] = 0;
   assign ecchmatrix[3][77] = 0;
   assign ecchmatrix[4][77] = 1;
   assign ecchmatrix[5][77] = 0;
   assign ecchmatrix[6][77] = 1;
   assign ecchmatrix[7][77] = 1;
   assign ecchmatrix[8][77] = 0;
   assign ecchmatrix[0][78] = 0;
   assign ecchmatrix[1][78] = 0;
   assign ecchmatrix[2][78] = 0;
   assign ecchmatrix[3][78] = 0;
   assign ecchmatrix[4][78] = 1;
   assign ecchmatrix[5][78] = 0;
   assign ecchmatrix[6][78] = 1;
   assign ecchmatrix[7][78] = 0;
   assign ecchmatrix[8][78] = 1;
   assign ecchmatrix[0][79] = 0;
   assign ecchmatrix[1][79] = 0;
   assign ecchmatrix[2][79] = 0;
   assign ecchmatrix[3][79] = 0;
   assign ecchmatrix[4][79] = 1;
   assign ecchmatrix[5][79] = 0;
   assign ecchmatrix[6][79] = 0;
   assign ecchmatrix[7][79] = 1;
   assign ecchmatrix[8][79] = 1;
   assign ecchmatrix[0][80] = 0;
   assign ecchmatrix[1][80] = 0;
   assign ecchmatrix[2][80] = 0;
   assign ecchmatrix[3][80] = 0;
   assign ecchmatrix[4][80] = 0;
   assign ecchmatrix[5][80] = 1;
   assign ecchmatrix[6][80] = 1;
   assign ecchmatrix[7][80] = 1;
   assign ecchmatrix[8][80] = 0;
   assign ecchmatrix[0][81] = 0;
   assign ecchmatrix[1][81] = 0;
   assign ecchmatrix[2][81] = 0;
   assign ecchmatrix[3][81] = 0;
   assign ecchmatrix[4][81] = 0;
   assign ecchmatrix[5][81] = 1;
   assign ecchmatrix[6][81] = 1;
   assign ecchmatrix[7][81] = 0;
   assign ecchmatrix[8][81] = 1;
   assign ecchmatrix[0][82] = 0;
   assign ecchmatrix[1][82] = 0;
   assign ecchmatrix[2][82] = 0;
   assign ecchmatrix[3][82] = 0;
   assign ecchmatrix[4][82] = 0;
   assign ecchmatrix[5][82] = 1;
   assign ecchmatrix[6][82] = 0;
   assign ecchmatrix[7][82] = 1;
   assign ecchmatrix[8][82] = 1;
   assign ecchmatrix[0][83] = 0;
   assign ecchmatrix[1][83] = 0;
   assign ecchmatrix[2][83] = 0;
   assign ecchmatrix[3][83] = 0;
   assign ecchmatrix[4][83] = 0;
   assign ecchmatrix[5][83] = 0;
   assign ecchmatrix[6][83] = 1;
   assign ecchmatrix[7][83] = 1;
   assign ecchmatrix[8][83] = 1;
   assign ecchmatrix[0][84] = 1;
   assign ecchmatrix[1][84] = 1;
   assign ecchmatrix[2][84] = 1;
   assign ecchmatrix[3][84] = 1;
   assign ecchmatrix[4][84] = 1;
   assign ecchmatrix[5][84] = 0;
   assign ecchmatrix[6][84] = 0;
   assign ecchmatrix[7][84] = 0;
   assign ecchmatrix[8][84] = 0;
   assign ecchmatrix[0][85] = 1;
   assign ecchmatrix[1][85] = 1;
   assign ecchmatrix[2][85] = 1;
   assign ecchmatrix[3][85] = 1;
   assign ecchmatrix[4][85] = 0;
   assign ecchmatrix[5][85] = 1;
   assign ecchmatrix[6][85] = 0;
   assign ecchmatrix[7][85] = 0;
   assign ecchmatrix[8][85] = 0;
   assign ecchmatrix[0][86] = 1;
   assign ecchmatrix[1][86] = 1;
   assign ecchmatrix[2][86] = 1;
   assign ecchmatrix[3][86] = 1;
   assign ecchmatrix[4][86] = 0;
   assign ecchmatrix[5][86] = 0;
   assign ecchmatrix[6][86] = 1;
   assign ecchmatrix[7][86] = 0;
   assign ecchmatrix[8][86] = 0;
   assign ecchmatrix[0][87] = 1;
   assign ecchmatrix[1][87] = 1;
   assign ecchmatrix[2][87] = 1;
   assign ecchmatrix[3][87] = 1;
   assign ecchmatrix[4][87] = 0;
   assign ecchmatrix[5][87] = 0;
   assign ecchmatrix[6][87] = 0;
   assign ecchmatrix[7][87] = 1;
   assign ecchmatrix[8][87] = 0;
   assign ecchmatrix[0][88] = 1;
   assign ecchmatrix[1][88] = 1;
   assign ecchmatrix[2][88] = 1;
   assign ecchmatrix[3][88] = 1;
   assign ecchmatrix[4][88] = 0;
   assign ecchmatrix[5][88] = 0;
   assign ecchmatrix[6][88] = 0;
   assign ecchmatrix[7][88] = 0;
   assign ecchmatrix[8][88] = 1;
   assign ecchmatrix[0][89] = 1;
   assign ecchmatrix[1][89] = 1;
   assign ecchmatrix[2][89] = 1;
   assign ecchmatrix[3][89] = 0;
   assign ecchmatrix[4][89] = 1;
   assign ecchmatrix[5][89] = 1;
   assign ecchmatrix[6][89] = 0;
   assign ecchmatrix[7][89] = 0;
   assign ecchmatrix[8][89] = 0;
   assign ecchmatrix[0][90] = 1;
   assign ecchmatrix[1][90] = 1;
   assign ecchmatrix[2][90] = 1;
   assign ecchmatrix[3][90] = 0;
   assign ecchmatrix[4][90] = 1;
   assign ecchmatrix[5][90] = 0;
   assign ecchmatrix[6][90] = 1;
   assign ecchmatrix[7][90] = 0;
   assign ecchmatrix[8][90] = 0;
   assign ecchmatrix[0][91] = 1;
   assign ecchmatrix[1][91] = 1;
   assign ecchmatrix[2][91] = 1;
   assign ecchmatrix[3][91] = 0;
   assign ecchmatrix[4][91] = 1;
   assign ecchmatrix[5][91] = 0;
   assign ecchmatrix[6][91] = 0;
   assign ecchmatrix[7][91] = 1;
   assign ecchmatrix[8][91] = 0;
   assign ecchmatrix[0][92] = 1;
   assign ecchmatrix[1][92] = 1;
   assign ecchmatrix[2][92] = 1;
   assign ecchmatrix[3][92] = 0;
   assign ecchmatrix[4][92] = 1;
   assign ecchmatrix[5][92] = 0;
   assign ecchmatrix[6][92] = 0;
   assign ecchmatrix[7][92] = 0;
   assign ecchmatrix[8][92] = 1;
   assign ecchmatrix[0][93] = 1;
   assign ecchmatrix[1][93] = 1;
   assign ecchmatrix[2][93] = 1;
   assign ecchmatrix[3][93] = 0;
   assign ecchmatrix[4][93] = 0;
   assign ecchmatrix[5][93] = 1;
   assign ecchmatrix[6][93] = 1;
   assign ecchmatrix[7][93] = 0;
   assign ecchmatrix[8][93] = 0;
   assign ecchmatrix[0][94] = 1;
   assign ecchmatrix[1][94] = 1;
   assign ecchmatrix[2][94] = 1;
   assign ecchmatrix[3][94] = 0;
   assign ecchmatrix[4][94] = 0;
   assign ecchmatrix[5][94] = 1;
   assign ecchmatrix[6][94] = 0;
   assign ecchmatrix[7][94] = 1;
   assign ecchmatrix[8][94] = 0;
   assign ecchmatrix[0][95] = 1;
   assign ecchmatrix[1][95] = 1;
   assign ecchmatrix[2][95] = 1;
   assign ecchmatrix[3][95] = 0;
   assign ecchmatrix[4][95] = 0;
   assign ecchmatrix[5][95] = 1;
   assign ecchmatrix[6][95] = 0;
   assign ecchmatrix[7][95] = 0;
   assign ecchmatrix[8][95] = 1;
   assign ecchmatrix[0][96] = 1;
   assign ecchmatrix[1][96] = 1;
   assign ecchmatrix[2][96] = 1;
   assign ecchmatrix[3][96] = 0;
   assign ecchmatrix[4][96] = 0;
   assign ecchmatrix[5][96] = 0;
   assign ecchmatrix[6][96] = 1;
   assign ecchmatrix[7][96] = 1;
   assign ecchmatrix[8][96] = 0;
   assign ecchmatrix[0][97] = 1;
   assign ecchmatrix[1][97] = 1;
   assign ecchmatrix[2][97] = 1;
   assign ecchmatrix[3][97] = 0;
   assign ecchmatrix[4][97] = 0;
   assign ecchmatrix[5][97] = 0;
   assign ecchmatrix[6][97] = 1;
   assign ecchmatrix[7][97] = 0;
   assign ecchmatrix[8][97] = 1;
   assign ecchmatrix[0][98] = 1;
   assign ecchmatrix[1][98] = 1;
   assign ecchmatrix[2][98] = 1;
   assign ecchmatrix[3][98] = 0;
   assign ecchmatrix[4][98] = 0;
   assign ecchmatrix[5][98] = 0;
   assign ecchmatrix[6][98] = 0;
   assign ecchmatrix[7][98] = 1;
   assign ecchmatrix[8][98] = 1;
   assign ecchmatrix[0][99] = 1;
   assign ecchmatrix[1][99] = 1;
   assign ecchmatrix[2][99] = 0;
   assign ecchmatrix[3][99] = 1;
   assign ecchmatrix[4][99] = 1;
   assign ecchmatrix[5][99] = 1;
   assign ecchmatrix[6][99] = 0;
   assign ecchmatrix[7][99] = 0;
   assign ecchmatrix[8][99] = 0;
   assign ecchmatrix[0][100] = 1;
   assign ecchmatrix[1][100] = 1;
   assign ecchmatrix[2][100] = 0;
   assign ecchmatrix[3][100] = 1;
   assign ecchmatrix[4][100] = 1;
   assign ecchmatrix[5][100] = 0;
   assign ecchmatrix[6][100] = 1;
   assign ecchmatrix[7][100] = 0;
   assign ecchmatrix[8][100] = 0;
   assign ecchmatrix[0][101] = 1;
   assign ecchmatrix[1][101] = 1;
   assign ecchmatrix[2][101] = 0;
   assign ecchmatrix[3][101] = 1;
   assign ecchmatrix[4][101] = 1;
   assign ecchmatrix[5][101] = 0;
   assign ecchmatrix[6][101] = 0;
   assign ecchmatrix[7][101] = 1;
   assign ecchmatrix[8][101] = 0;
   assign ecchmatrix[0][102] = 1;
   assign ecchmatrix[1][102] = 1;
   assign ecchmatrix[2][102] = 0;
   assign ecchmatrix[3][102] = 1;
   assign ecchmatrix[4][102] = 1;
   assign ecchmatrix[5][102] = 0;
   assign ecchmatrix[6][102] = 0;
   assign ecchmatrix[7][102] = 0;
   assign ecchmatrix[8][102] = 1;
   assign ecchmatrix[0][103] = 1;
   assign ecchmatrix[1][103] = 1;
   assign ecchmatrix[2][103] = 0;
   assign ecchmatrix[3][103] = 1;
   assign ecchmatrix[4][103] = 0;
   assign ecchmatrix[5][103] = 1;
   assign ecchmatrix[6][103] = 1;
   assign ecchmatrix[7][103] = 0;
   assign ecchmatrix[8][103] = 0;
   assign ecchmatrix[0][104] = 1;
   assign ecchmatrix[1][104] = 1;
   assign ecchmatrix[2][104] = 0;
   assign ecchmatrix[3][104] = 1;
   assign ecchmatrix[4][104] = 0;
   assign ecchmatrix[5][104] = 1;
   assign ecchmatrix[6][104] = 0;
   assign ecchmatrix[7][104] = 1;
   assign ecchmatrix[8][104] = 0;
   assign ecchmatrix[0][105] = 1;
   assign ecchmatrix[1][105] = 1;
   assign ecchmatrix[2][105] = 0;
   assign ecchmatrix[3][105] = 1;
   assign ecchmatrix[4][105] = 0;
   assign ecchmatrix[5][105] = 1;
   assign ecchmatrix[6][105] = 0;
   assign ecchmatrix[7][105] = 0;
   assign ecchmatrix[8][105] = 1;
   assign ecchmatrix[0][106] = 1;
   assign ecchmatrix[1][106] = 1;
   assign ecchmatrix[2][106] = 0;
   assign ecchmatrix[3][106] = 1;
   assign ecchmatrix[4][106] = 0;
   assign ecchmatrix[5][106] = 0;
   assign ecchmatrix[6][106] = 1;
   assign ecchmatrix[7][106] = 1;
   assign ecchmatrix[8][106] = 0;
   assign ecchmatrix[0][107] = 1;
   assign ecchmatrix[1][107] = 1;
   assign ecchmatrix[2][107] = 0;
   assign ecchmatrix[3][107] = 1;
   assign ecchmatrix[4][107] = 0;
   assign ecchmatrix[5][107] = 0;
   assign ecchmatrix[6][107] = 1;
   assign ecchmatrix[7][107] = 0;
   assign ecchmatrix[8][107] = 1;
   assign ecchmatrix[0][108] = 1;
   assign ecchmatrix[1][108] = 1;
   assign ecchmatrix[2][108] = 0;
   assign ecchmatrix[3][108] = 1;
   assign ecchmatrix[4][108] = 0;
   assign ecchmatrix[5][108] = 0;
   assign ecchmatrix[6][108] = 0;
   assign ecchmatrix[7][108] = 1;
   assign ecchmatrix[8][108] = 1;
   assign ecchmatrix[0][109] = 1;
   assign ecchmatrix[1][109] = 1;
   assign ecchmatrix[2][109] = 0;
   assign ecchmatrix[3][109] = 0;
   assign ecchmatrix[4][109] = 1;
   assign ecchmatrix[5][109] = 1;
   assign ecchmatrix[6][109] = 1;
   assign ecchmatrix[7][109] = 0;
   assign ecchmatrix[8][109] = 0;
   assign ecchmatrix[0][110] = 1;
   assign ecchmatrix[1][110] = 1;
   assign ecchmatrix[2][110] = 0;
   assign ecchmatrix[3][110] = 0;
   assign ecchmatrix[4][110] = 1;
   assign ecchmatrix[5][110] = 1;
   assign ecchmatrix[6][110] = 0;
   assign ecchmatrix[7][110] = 1;
   assign ecchmatrix[8][110] = 0;
   assign ecchmatrix[0][111] = 1;
   assign ecchmatrix[1][111] = 1;
   assign ecchmatrix[2][111] = 0;
   assign ecchmatrix[3][111] = 0;
   assign ecchmatrix[4][111] = 1;
   assign ecchmatrix[5][111] = 1;
   assign ecchmatrix[6][111] = 0;
   assign ecchmatrix[7][111] = 0;
   assign ecchmatrix[8][111] = 1;
   assign ecchmatrix[0][112] = 1;
   assign ecchmatrix[1][112] = 1;
   assign ecchmatrix[2][112] = 0;
   assign ecchmatrix[3][112] = 0;
   assign ecchmatrix[4][112] = 1;
   assign ecchmatrix[5][112] = 0;
   assign ecchmatrix[6][112] = 1;
   assign ecchmatrix[7][112] = 1;
   assign ecchmatrix[8][112] = 0;
   assign ecchmatrix[0][113] = 1;
   assign ecchmatrix[1][113] = 1;
   assign ecchmatrix[2][113] = 0;
   assign ecchmatrix[3][113] = 0;
   assign ecchmatrix[4][113] = 1;
   assign ecchmatrix[5][113] = 0;
   assign ecchmatrix[6][113] = 1;
   assign ecchmatrix[7][113] = 0;
   assign ecchmatrix[8][113] = 1;
   assign ecchmatrix[0][114] = 1;
   assign ecchmatrix[1][114] = 1;
   assign ecchmatrix[2][114] = 0;
   assign ecchmatrix[3][114] = 0;
   assign ecchmatrix[4][114] = 1;
   assign ecchmatrix[5][114] = 0;
   assign ecchmatrix[6][114] = 0;
   assign ecchmatrix[7][114] = 1;
   assign ecchmatrix[8][114] = 1;
   assign ecchmatrix[0][115] = 1;
   assign ecchmatrix[1][115] = 1;
   assign ecchmatrix[2][115] = 0;
   assign ecchmatrix[3][115] = 0;
   assign ecchmatrix[4][115] = 0;
   assign ecchmatrix[5][115] = 1;
   assign ecchmatrix[6][115] = 1;
   assign ecchmatrix[7][115] = 1;
   assign ecchmatrix[8][115] = 0;
   assign ecchmatrix[0][116] = 1;
   assign ecchmatrix[1][116] = 1;
   assign ecchmatrix[2][116] = 0;
   assign ecchmatrix[3][116] = 0;
   assign ecchmatrix[4][116] = 0;
   assign ecchmatrix[5][116] = 1;
   assign ecchmatrix[6][116] = 1;
   assign ecchmatrix[7][116] = 0;
   assign ecchmatrix[8][116] = 1;
   assign ecchmatrix[0][117] = 1;
   assign ecchmatrix[1][117] = 1;
   assign ecchmatrix[2][117] = 0;
   assign ecchmatrix[3][117] = 0;
   assign ecchmatrix[4][117] = 0;
   assign ecchmatrix[5][117] = 1;
   assign ecchmatrix[6][117] = 0;
   assign ecchmatrix[7][117] = 1;
   assign ecchmatrix[8][117] = 1;
   assign ecchmatrix[0][118] = 1;
   assign ecchmatrix[1][118] = 1;
   assign ecchmatrix[2][118] = 0;
   assign ecchmatrix[3][118] = 0;
   assign ecchmatrix[4][118] = 0;
   assign ecchmatrix[5][118] = 0;
   assign ecchmatrix[6][118] = 1;
   assign ecchmatrix[7][118] = 1;
   assign ecchmatrix[8][118] = 1;
   assign ecchmatrix[0][119] = 1;
   assign ecchmatrix[1][119] = 0;
   assign ecchmatrix[2][119] = 1;
   assign ecchmatrix[3][119] = 1;
   assign ecchmatrix[4][119] = 1;
   assign ecchmatrix[5][119] = 1;
   assign ecchmatrix[6][119] = 0;
   assign ecchmatrix[7][119] = 0;
   assign ecchmatrix[8][119] = 0;
   assign ecchmatrix[0][120] = 1;
   assign ecchmatrix[1][120] = 0;
   assign ecchmatrix[2][120] = 1;
   assign ecchmatrix[3][120] = 1;
   assign ecchmatrix[4][120] = 1;
   assign ecchmatrix[5][120] = 0;
   assign ecchmatrix[6][120] = 1;
   assign ecchmatrix[7][120] = 0;
   assign ecchmatrix[8][120] = 0;
   assign ecchmatrix[0][121] = 1;
   assign ecchmatrix[1][121] = 0;
   assign ecchmatrix[2][121] = 1;
   assign ecchmatrix[3][121] = 1;
   assign ecchmatrix[4][121] = 1;
   assign ecchmatrix[5][121] = 0;
   assign ecchmatrix[6][121] = 0;
   assign ecchmatrix[7][121] = 1;
   assign ecchmatrix[8][121] = 0;
   assign ecchmatrix[0][122] = 1;
   assign ecchmatrix[1][122] = 0;
   assign ecchmatrix[2][122] = 1;
   assign ecchmatrix[3][122] = 1;
   assign ecchmatrix[4][122] = 1;
   assign ecchmatrix[5][122] = 0;
   assign ecchmatrix[6][122] = 0;
   assign ecchmatrix[7][122] = 0;
   assign ecchmatrix[8][122] = 1;
   assign ecchmatrix[0][123] = 1;
   assign ecchmatrix[1][123] = 0;
   assign ecchmatrix[2][123] = 1;
   assign ecchmatrix[3][123] = 1;
   assign ecchmatrix[4][123] = 0;
   assign ecchmatrix[5][123] = 1;
   assign ecchmatrix[6][123] = 1;
   assign ecchmatrix[7][123] = 0;
   assign ecchmatrix[8][123] = 0;
   assign ecchmatrix[0][124] = 1;
   assign ecchmatrix[1][124] = 0;
   assign ecchmatrix[2][124] = 1;
   assign ecchmatrix[3][124] = 1;
   assign ecchmatrix[4][124] = 0;
   assign ecchmatrix[5][124] = 1;
   assign ecchmatrix[6][124] = 0;
   assign ecchmatrix[7][124] = 1;
   assign ecchmatrix[8][124] = 0;
   assign ecchmatrix[0][125] = 1;
   assign ecchmatrix[1][125] = 0;
   assign ecchmatrix[2][125] = 1;
   assign ecchmatrix[3][125] = 1;
   assign ecchmatrix[4][125] = 0;
   assign ecchmatrix[5][125] = 1;
   assign ecchmatrix[6][125] = 0;
   assign ecchmatrix[7][125] = 0;
   assign ecchmatrix[8][125] = 1;
   assign ecchmatrix[0][126] = 1;
   assign ecchmatrix[1][126] = 0;
   assign ecchmatrix[2][126] = 1;
   assign ecchmatrix[3][126] = 1;
   assign ecchmatrix[4][126] = 0;
   assign ecchmatrix[5][126] = 0;
   assign ecchmatrix[6][126] = 1;
   assign ecchmatrix[7][126] = 1;
   assign ecchmatrix[8][126] = 0;
   assign ecchmatrix[0][127] = 1;
   assign ecchmatrix[1][127] = 0;
   assign ecchmatrix[2][127] = 1;
   assign ecchmatrix[3][127] = 1;
   assign ecchmatrix[4][127] = 0;
   assign ecchmatrix[5][127] = 0;
   assign ecchmatrix[6][127] = 1;
   assign ecchmatrix[7][127] = 0;
   assign ecchmatrix[8][127] = 1;
   assign ecchmatrix[0][128] = 1;
   assign ecchmatrix[1][128] = 0;
   assign ecchmatrix[2][128] = 1;
   assign ecchmatrix[3][128] = 1;
   assign ecchmatrix[4][128] = 0;
   assign ecchmatrix[5][128] = 0;
   assign ecchmatrix[6][128] = 0;
   assign ecchmatrix[7][128] = 1;
   assign ecchmatrix[8][128] = 1;
   assign ecchmatrix[0][129] = 1;
   assign ecchmatrix[1][129] = 0;
   assign ecchmatrix[2][129] = 1;
   assign ecchmatrix[3][129] = 0;
   assign ecchmatrix[4][129] = 1;
   assign ecchmatrix[5][129] = 1;
   assign ecchmatrix[6][129] = 1;
   assign ecchmatrix[7][129] = 0;
   assign ecchmatrix[8][129] = 0;
   assign ecchmatrix[0][130] = 1;
   assign ecchmatrix[1][130] = 0;
   assign ecchmatrix[2][130] = 1;
   assign ecchmatrix[3][130] = 0;
   assign ecchmatrix[4][130] = 1;
   assign ecchmatrix[5][130] = 1;
   assign ecchmatrix[6][130] = 0;
   assign ecchmatrix[7][130] = 1;
   assign ecchmatrix[8][130] = 0;
   assign ecchmatrix[0][131] = 1;
   assign ecchmatrix[1][131] = 0;
   assign ecchmatrix[2][131] = 1;
   assign ecchmatrix[3][131] = 0;
   assign ecchmatrix[4][131] = 1;
   assign ecchmatrix[5][131] = 1;
   assign ecchmatrix[6][131] = 0;
   assign ecchmatrix[7][131] = 0;
   assign ecchmatrix[8][131] = 1;
   assign ecchmatrix[0][132] = 1;
   assign ecchmatrix[1][132] = 0;
   assign ecchmatrix[2][132] = 1;
   assign ecchmatrix[3][132] = 0;
   assign ecchmatrix[4][132] = 1;
   assign ecchmatrix[5][132] = 0;
   assign ecchmatrix[6][132] = 1;
   assign ecchmatrix[7][132] = 1;
   assign ecchmatrix[8][132] = 0;
   assign ecchmatrix[0][133] = 1;
   assign ecchmatrix[1][133] = 0;
   assign ecchmatrix[2][133] = 1;
   assign ecchmatrix[3][133] = 0;
   assign ecchmatrix[4][133] = 1;
   assign ecchmatrix[5][133] = 0;
   assign ecchmatrix[6][133] = 1;
   assign ecchmatrix[7][133] = 0;
   assign ecchmatrix[8][133] = 1;
   assign ecchmatrix[0][134] = 1;
   assign ecchmatrix[1][134] = 0;
   assign ecchmatrix[2][134] = 1;
   assign ecchmatrix[3][134] = 0;
   assign ecchmatrix[4][134] = 1;
   assign ecchmatrix[5][134] = 0;
   assign ecchmatrix[6][134] = 0;
   assign ecchmatrix[7][134] = 1;
   assign ecchmatrix[8][134] = 1;
   assign ecchmatrix[0][135] = 1;
   assign ecchmatrix[1][135] = 0;
   assign ecchmatrix[2][135] = 1;
   assign ecchmatrix[3][135] = 0;
   assign ecchmatrix[4][135] = 0;
   assign ecchmatrix[5][135] = 1;
   assign ecchmatrix[6][135] = 1;
   assign ecchmatrix[7][135] = 1;
   assign ecchmatrix[8][135] = 0;
   assign ecchmatrix[0][136] = 1;
   assign ecchmatrix[1][136] = 0;
   assign ecchmatrix[2][136] = 1;
   assign ecchmatrix[3][136] = 0;
   assign ecchmatrix[4][136] = 0;
   assign ecchmatrix[5][136] = 1;
   assign ecchmatrix[6][136] = 1;
   assign ecchmatrix[7][136] = 0;
   assign ecchmatrix[8][136] = 1;
   assign ecchmatrix[0][137] = 1;
   assign ecchmatrix[1][137] = 0;
   assign ecchmatrix[2][137] = 1;
   assign ecchmatrix[3][137] = 0;
   assign ecchmatrix[4][137] = 0;
   assign ecchmatrix[5][137] = 1;
   assign ecchmatrix[6][137] = 0;
   assign ecchmatrix[7][137] = 1;
   assign ecchmatrix[8][137] = 1;
   assign ecchmatrix[0][138] = 1;
   assign ecchmatrix[1][138] = 0;
   assign ecchmatrix[2][138] = 1;
   assign ecchmatrix[3][138] = 0;
   assign ecchmatrix[4][138] = 0;
   assign ecchmatrix[5][138] = 0;
   assign ecchmatrix[6][138] = 1;
   assign ecchmatrix[7][138] = 1;
   assign ecchmatrix[8][138] = 1;
   assign ecchmatrix[0][139] = 1;
   assign ecchmatrix[1][139] = 0;
   assign ecchmatrix[2][139] = 0;
   assign ecchmatrix[3][139] = 1;
   assign ecchmatrix[4][139] = 1;
   assign ecchmatrix[5][139] = 1;
   assign ecchmatrix[6][139] = 1;
   assign ecchmatrix[7][139] = 0;
   assign ecchmatrix[8][139] = 0;
   assign ecchmatrix[0][140] = 1;
   assign ecchmatrix[1][140] = 0;
   assign ecchmatrix[2][140] = 0;
   assign ecchmatrix[3][140] = 1;
   assign ecchmatrix[4][140] = 1;
   assign ecchmatrix[5][140] = 1;
   assign ecchmatrix[6][140] = 0;
   assign ecchmatrix[7][140] = 1;
   assign ecchmatrix[8][140] = 0;
   assign ecchmatrix[0][141] = 1;
   assign ecchmatrix[1][141] = 0;
   assign ecchmatrix[2][141] = 0;
   assign ecchmatrix[3][141] = 1;
   assign ecchmatrix[4][141] = 1;
   assign ecchmatrix[5][141] = 1;
   assign ecchmatrix[6][141] = 0;
   assign ecchmatrix[7][141] = 0;
   assign ecchmatrix[8][141] = 1;
   assign ecchmatrix[0][142] = 1;
   assign ecchmatrix[1][142] = 0;
   assign ecchmatrix[2][142] = 0;
   assign ecchmatrix[3][142] = 1;
   assign ecchmatrix[4][142] = 1;
   assign ecchmatrix[5][142] = 0;
   assign ecchmatrix[6][142] = 1;
   assign ecchmatrix[7][142] = 1;
   assign ecchmatrix[8][142] = 0;
   assign ecchmatrix[0][143] = 1;
   assign ecchmatrix[1][143] = 0;
   assign ecchmatrix[2][143] = 0;
   assign ecchmatrix[3][143] = 1;
   assign ecchmatrix[4][143] = 1;
   assign ecchmatrix[5][143] = 0;
   assign ecchmatrix[6][143] = 1;
   assign ecchmatrix[7][143] = 0;
   assign ecchmatrix[8][143] = 1;
   assign ecchmatrix[0][144] = 1;
   assign ecchmatrix[1][144] = 0;
   assign ecchmatrix[2][144] = 0;
   assign ecchmatrix[3][144] = 1;
   assign ecchmatrix[4][144] = 1;
   assign ecchmatrix[5][144] = 0;
   assign ecchmatrix[6][144] = 0;
   assign ecchmatrix[7][144] = 1;
   assign ecchmatrix[8][144] = 1;
   assign ecchmatrix[0][145] = 1;
   assign ecchmatrix[1][145] = 0;
   assign ecchmatrix[2][145] = 0;
   assign ecchmatrix[3][145] = 1;
   assign ecchmatrix[4][145] = 0;
   assign ecchmatrix[5][145] = 1;
   assign ecchmatrix[6][145] = 1;
   assign ecchmatrix[7][145] = 1;
   assign ecchmatrix[8][145] = 0;
   assign ecchmatrix[0][146] = 1;
   assign ecchmatrix[1][146] = 0;
   assign ecchmatrix[2][146] = 0;
   assign ecchmatrix[3][146] = 1;
   assign ecchmatrix[4][146] = 0;
   assign ecchmatrix[5][146] = 1;
   assign ecchmatrix[6][146] = 1;
   assign ecchmatrix[7][146] = 0;
   assign ecchmatrix[8][146] = 1;
   assign ecchmatrix[0][147] = 1;
   assign ecchmatrix[1][147] = 0;
   assign ecchmatrix[2][147] = 0;
   assign ecchmatrix[3][147] = 1;
   assign ecchmatrix[4][147] = 0;
   assign ecchmatrix[5][147] = 1;
   assign ecchmatrix[6][147] = 0;
   assign ecchmatrix[7][147] = 1;
   assign ecchmatrix[8][147] = 1;
   assign ecchmatrix[0][148] = 1;
   assign ecchmatrix[1][148] = 0;
   assign ecchmatrix[2][148] = 0;
   assign ecchmatrix[3][148] = 1;
   assign ecchmatrix[4][148] = 0;
   assign ecchmatrix[5][148] = 0;
   assign ecchmatrix[6][148] = 1;
   assign ecchmatrix[7][148] = 1;
   assign ecchmatrix[8][148] = 1;
   assign ecchmatrix[0][149] = 1;
   assign ecchmatrix[1][149] = 0;
   assign ecchmatrix[2][149] = 0;
   assign ecchmatrix[3][149] = 0;
   assign ecchmatrix[4][149] = 1;
   assign ecchmatrix[5][149] = 1;
   assign ecchmatrix[6][149] = 1;
   assign ecchmatrix[7][149] = 1;
   assign ecchmatrix[8][149] = 0;
   assign ecchmatrix[0][150] = 1;
   assign ecchmatrix[1][150] = 0;
   assign ecchmatrix[2][150] = 0;
   assign ecchmatrix[3][150] = 0;
   assign ecchmatrix[4][150] = 1;
   assign ecchmatrix[5][150] = 1;
   assign ecchmatrix[6][150] = 1;
   assign ecchmatrix[7][150] = 0;
   assign ecchmatrix[8][150] = 1;
   assign ecchmatrix[0][151] = 1;
   assign ecchmatrix[1][151] = 0;
   assign ecchmatrix[2][151] = 0;
   assign ecchmatrix[3][151] = 0;
   assign ecchmatrix[4][151] = 1;
   assign ecchmatrix[5][151] = 1;
   assign ecchmatrix[6][151] = 0;
   assign ecchmatrix[7][151] = 1;
   assign ecchmatrix[8][151] = 1;
   assign ecchmatrix[0][152] = 1;
   assign ecchmatrix[1][152] = 0;
   assign ecchmatrix[2][152] = 0;
   assign ecchmatrix[3][152] = 0;
   assign ecchmatrix[4][152] = 1;
   assign ecchmatrix[5][152] = 0;
   assign ecchmatrix[6][152] = 1;
   assign ecchmatrix[7][152] = 1;
   assign ecchmatrix[8][152] = 1;
   assign ecchmatrix[0][153] = 1;
   assign ecchmatrix[1][153] = 0;
   assign ecchmatrix[2][153] = 0;
   assign ecchmatrix[3][153] = 0;
   assign ecchmatrix[4][153] = 0;
   assign ecchmatrix[5][153] = 1;
   assign ecchmatrix[6][153] = 1;
   assign ecchmatrix[7][153] = 1;
   assign ecchmatrix[8][153] = 1;
   assign ecchmatrix[0][154] = 0;
   assign ecchmatrix[1][154] = 1;
   assign ecchmatrix[2][154] = 1;
   assign ecchmatrix[3][154] = 1;
   assign ecchmatrix[4][154] = 1;
   assign ecchmatrix[5][154] = 1;
   assign ecchmatrix[6][154] = 0;
   assign ecchmatrix[7][154] = 0;
   assign ecchmatrix[8][154] = 0;
   assign ecchmatrix[0][155] = 0;
   assign ecchmatrix[1][155] = 1;
   assign ecchmatrix[2][155] = 1;
   assign ecchmatrix[3][155] = 1;
   assign ecchmatrix[4][155] = 1;
   assign ecchmatrix[5][155] = 0;
   assign ecchmatrix[6][155] = 1;
   assign ecchmatrix[7][155] = 0;
   assign ecchmatrix[8][155] = 0;
   assign ecchmatrix[0][156] = 0;
   assign ecchmatrix[1][156] = 1;
   assign ecchmatrix[2][156] = 1;
   assign ecchmatrix[3][156] = 1;
   assign ecchmatrix[4][156] = 1;
   assign ecchmatrix[5][156] = 0;
   assign ecchmatrix[6][156] = 0;
   assign ecchmatrix[7][156] = 1;
   assign ecchmatrix[8][156] = 0;
   assign ecchmatrix[0][157] = 0;
   assign ecchmatrix[1][157] = 1;
   assign ecchmatrix[2][157] = 1;
   assign ecchmatrix[3][157] = 1;
   assign ecchmatrix[4][157] = 1;
   assign ecchmatrix[5][157] = 0;
   assign ecchmatrix[6][157] = 0;
   assign ecchmatrix[7][157] = 0;
   assign ecchmatrix[8][157] = 1;
   assign ecchmatrix[0][158] = 0;
   assign ecchmatrix[1][158] = 1;
   assign ecchmatrix[2][158] = 1;
   assign ecchmatrix[3][158] = 1;
   assign ecchmatrix[4][158] = 0;
   assign ecchmatrix[5][158] = 1;
   assign ecchmatrix[6][158] = 1;
   assign ecchmatrix[7][158] = 0;
   assign ecchmatrix[8][158] = 0;
   assign ecchmatrix[0][159] = 0;
   assign ecchmatrix[1][159] = 1;
   assign ecchmatrix[2][159] = 1;
   assign ecchmatrix[3][159] = 1;
   assign ecchmatrix[4][159] = 0;
   assign ecchmatrix[5][159] = 1;
   assign ecchmatrix[6][159] = 0;
   assign ecchmatrix[7][159] = 1;
   assign ecchmatrix[8][159] = 0;
   assign ecchmatrix[0][160] = 0;
   assign ecchmatrix[1][160] = 1;
   assign ecchmatrix[2][160] = 1;
   assign ecchmatrix[3][160] = 1;
   assign ecchmatrix[4][160] = 0;
   assign ecchmatrix[5][160] = 1;
   assign ecchmatrix[6][160] = 0;
   assign ecchmatrix[7][160] = 0;
   assign ecchmatrix[8][160] = 1;
   assign ecchmatrix[0][161] = 0;
   assign ecchmatrix[1][161] = 1;
   assign ecchmatrix[2][161] = 1;
   assign ecchmatrix[3][161] = 1;
   assign ecchmatrix[4][161] = 0;
   assign ecchmatrix[5][161] = 0;
   assign ecchmatrix[6][161] = 1;
   assign ecchmatrix[7][161] = 1;
   assign ecchmatrix[8][161] = 0;
   assign ecchmatrix[0][162] = 0;
   assign ecchmatrix[1][162] = 1;
   assign ecchmatrix[2][162] = 1;
   assign ecchmatrix[3][162] = 1;
   assign ecchmatrix[4][162] = 0;
   assign ecchmatrix[5][162] = 0;
   assign ecchmatrix[6][162] = 1;
   assign ecchmatrix[7][162] = 0;
   assign ecchmatrix[8][162] = 1;
   assign ecchmatrix[0][163] = 0;
   assign ecchmatrix[1][163] = 1;
   assign ecchmatrix[2][163] = 1;
   assign ecchmatrix[3][163] = 1;
   assign ecchmatrix[4][163] = 0;
   assign ecchmatrix[5][163] = 0;
   assign ecchmatrix[6][163] = 0;
   assign ecchmatrix[7][163] = 1;
   assign ecchmatrix[8][163] = 1;
   assign ecchmatrix[0][164] = 0;
   assign ecchmatrix[1][164] = 1;
   assign ecchmatrix[2][164] = 1;
   assign ecchmatrix[3][164] = 0;
   assign ecchmatrix[4][164] = 1;
   assign ecchmatrix[5][164] = 1;
   assign ecchmatrix[6][164] = 1;
   assign ecchmatrix[7][164] = 0;
   assign ecchmatrix[8][164] = 0;
   assign ecchmatrix[0][165] = 0;
   assign ecchmatrix[1][165] = 1;
   assign ecchmatrix[2][165] = 1;
   assign ecchmatrix[3][165] = 0;
   assign ecchmatrix[4][165] = 1;
   assign ecchmatrix[5][165] = 1;
   assign ecchmatrix[6][165] = 0;
   assign ecchmatrix[7][165] = 1;
   assign ecchmatrix[8][165] = 0;
   assign ecchmatrix[0][166] = 0;
   assign ecchmatrix[1][166] = 1;
   assign ecchmatrix[2][166] = 1;
   assign ecchmatrix[3][166] = 0;
   assign ecchmatrix[4][166] = 1;
   assign ecchmatrix[5][166] = 1;
   assign ecchmatrix[6][166] = 0;
   assign ecchmatrix[7][166] = 0;
   assign ecchmatrix[8][166] = 1;
   assign ecchmatrix[0][167] = 0;
   assign ecchmatrix[1][167] = 1;
   assign ecchmatrix[2][167] = 1;
   assign ecchmatrix[3][167] = 0;
   assign ecchmatrix[4][167] = 1;
   assign ecchmatrix[5][167] = 0;
   assign ecchmatrix[6][167] = 1;
   assign ecchmatrix[7][167] = 1;
   assign ecchmatrix[8][167] = 0;
   assign ecchmatrix[0][168] = 0;
   assign ecchmatrix[1][168] = 1;
   assign ecchmatrix[2][168] = 1;
   assign ecchmatrix[3][168] = 0;
   assign ecchmatrix[4][168] = 1;
   assign ecchmatrix[5][168] = 0;
   assign ecchmatrix[6][168] = 1;
   assign ecchmatrix[7][168] = 0;
   assign ecchmatrix[8][168] = 1;
   assign ecchmatrix[0][169] = 0;
   assign ecchmatrix[1][169] = 1;
   assign ecchmatrix[2][169] = 1;
   assign ecchmatrix[3][169] = 0;
   assign ecchmatrix[4][169] = 1;
   assign ecchmatrix[5][169] = 0;
   assign ecchmatrix[6][169] = 0;
   assign ecchmatrix[7][169] = 1;
   assign ecchmatrix[8][169] = 1;
   assign ecchmatrix[0][170] = 0;
   assign ecchmatrix[1][170] = 1;
   assign ecchmatrix[2][170] = 1;
   assign ecchmatrix[3][170] = 0;
   assign ecchmatrix[4][170] = 0;
   assign ecchmatrix[5][170] = 1;
   assign ecchmatrix[6][170] = 1;
   assign ecchmatrix[7][170] = 1;
   assign ecchmatrix[8][170] = 0;
   assign ecchmatrix[0][171] = 0;
   assign ecchmatrix[1][171] = 1;
   assign ecchmatrix[2][171] = 1;
   assign ecchmatrix[3][171] = 0;
   assign ecchmatrix[4][171] = 0;
   assign ecchmatrix[5][171] = 1;
   assign ecchmatrix[6][171] = 1;
   assign ecchmatrix[7][171] = 0;
   assign ecchmatrix[8][171] = 1;
   assign ecchmatrix[0][172] = 0;
   assign ecchmatrix[1][172] = 1;
   assign ecchmatrix[2][172] = 1;
   assign ecchmatrix[3][172] = 0;
   assign ecchmatrix[4][172] = 0;
   assign ecchmatrix[5][172] = 1;
   assign ecchmatrix[6][172] = 0;
   assign ecchmatrix[7][172] = 1;
   assign ecchmatrix[8][172] = 1;
   assign ecchmatrix[0][173] = 0;
   assign ecchmatrix[1][173] = 1;
   assign ecchmatrix[2][173] = 1;
   assign ecchmatrix[3][173] = 0;
   assign ecchmatrix[4][173] = 0;
   assign ecchmatrix[5][173] = 0;
   assign ecchmatrix[6][173] = 1;
   assign ecchmatrix[7][173] = 1;
   assign ecchmatrix[8][173] = 1;
   assign ecchmatrix[0][174] = 0;
   assign ecchmatrix[1][174] = 1;
   assign ecchmatrix[2][174] = 0;
   assign ecchmatrix[3][174] = 1;
   assign ecchmatrix[4][174] = 1;
   assign ecchmatrix[5][174] = 1;
   assign ecchmatrix[6][174] = 1;
   assign ecchmatrix[7][174] = 0;
   assign ecchmatrix[8][174] = 0;
   assign ecchmatrix[0][175] = 0;
   assign ecchmatrix[1][175] = 1;
   assign ecchmatrix[2][175] = 0;
   assign ecchmatrix[3][175] = 1;
   assign ecchmatrix[4][175] = 1;
   assign ecchmatrix[5][175] = 1;
   assign ecchmatrix[6][175] = 0;
   assign ecchmatrix[7][175] = 1;
   assign ecchmatrix[8][175] = 0;
   assign ecchmatrix[0][176] = 0;
   assign ecchmatrix[1][176] = 1;
   assign ecchmatrix[2][176] = 0;
   assign ecchmatrix[3][176] = 1;
   assign ecchmatrix[4][176] = 1;
   assign ecchmatrix[5][176] = 1;
   assign ecchmatrix[6][176] = 0;
   assign ecchmatrix[7][176] = 0;
   assign ecchmatrix[8][176] = 1;
   assign ecchmatrix[0][177] = 0;
   assign ecchmatrix[1][177] = 1;
   assign ecchmatrix[2][177] = 0;
   assign ecchmatrix[3][177] = 1;
   assign ecchmatrix[4][177] = 1;
   assign ecchmatrix[5][177] = 0;
   assign ecchmatrix[6][177] = 1;
   assign ecchmatrix[7][177] = 1;
   assign ecchmatrix[8][177] = 0;
   assign ecchmatrix[0][178] = 0;
   assign ecchmatrix[1][178] = 1;
   assign ecchmatrix[2][178] = 0;
   assign ecchmatrix[3][178] = 1;
   assign ecchmatrix[4][178] = 1;
   assign ecchmatrix[5][178] = 0;
   assign ecchmatrix[6][178] = 1;
   assign ecchmatrix[7][178] = 0;
   assign ecchmatrix[8][178] = 1;
   assign ecchmatrix[0][179] = 0;
   assign ecchmatrix[1][179] = 1;
   assign ecchmatrix[2][179] = 0;
   assign ecchmatrix[3][179] = 1;
   assign ecchmatrix[4][179] = 1;
   assign ecchmatrix[5][179] = 0;
   assign ecchmatrix[6][179] = 0;
   assign ecchmatrix[7][179] = 1;
   assign ecchmatrix[8][179] = 1;
   assign ecchmatrix[0][180] = 0;
   assign ecchmatrix[1][180] = 1;
   assign ecchmatrix[2][180] = 0;
   assign ecchmatrix[3][180] = 1;
   assign ecchmatrix[4][180] = 0;
   assign ecchmatrix[5][180] = 1;
   assign ecchmatrix[6][180] = 1;
   assign ecchmatrix[7][180] = 1;
   assign ecchmatrix[8][180] = 0;
   assign ecchmatrix[0][181] = 0;
   assign ecchmatrix[1][181] = 1;
   assign ecchmatrix[2][181] = 0;
   assign ecchmatrix[3][181] = 1;
   assign ecchmatrix[4][181] = 0;
   assign ecchmatrix[5][181] = 1;
   assign ecchmatrix[6][181] = 1;
   assign ecchmatrix[7][181] = 0;
   assign ecchmatrix[8][181] = 1;
   assign ecchmatrix[0][182] = 0;
   assign ecchmatrix[1][182] = 1;
   assign ecchmatrix[2][182] = 0;
   assign ecchmatrix[3][182] = 1;
   assign ecchmatrix[4][182] = 0;
   assign ecchmatrix[5][182] = 1;
   assign ecchmatrix[6][182] = 0;
   assign ecchmatrix[7][182] = 1;
   assign ecchmatrix[8][182] = 1;
   assign ecchmatrix[0][183] = 0;
   assign ecchmatrix[1][183] = 1;
   assign ecchmatrix[2][183] = 0;
   assign ecchmatrix[3][183] = 1;
   assign ecchmatrix[4][183] = 0;
   assign ecchmatrix[5][183] = 0;
   assign ecchmatrix[6][183] = 1;
   assign ecchmatrix[7][183] = 1;
   assign ecchmatrix[8][183] = 1;
   assign ecchmatrix[0][184] = 0;
   assign ecchmatrix[1][184] = 1;
   assign ecchmatrix[2][184] = 0;
   assign ecchmatrix[3][184] = 0;
   assign ecchmatrix[4][184] = 1;
   assign ecchmatrix[5][184] = 1;
   assign ecchmatrix[6][184] = 1;
   assign ecchmatrix[7][184] = 1;
   assign ecchmatrix[8][184] = 0;
   assign ecchmatrix[0][185] = 0;
   assign ecchmatrix[1][185] = 1;
   assign ecchmatrix[2][185] = 0;
   assign ecchmatrix[3][185] = 0;
   assign ecchmatrix[4][185] = 1;
   assign ecchmatrix[5][185] = 1;
   assign ecchmatrix[6][185] = 1;
   assign ecchmatrix[7][185] = 0;
   assign ecchmatrix[8][185] = 1;
   assign ecchmatrix[0][186] = 0;
   assign ecchmatrix[1][186] = 1;
   assign ecchmatrix[2][186] = 0;
   assign ecchmatrix[3][186] = 0;
   assign ecchmatrix[4][186] = 1;
   assign ecchmatrix[5][186] = 1;
   assign ecchmatrix[6][186] = 0;
   assign ecchmatrix[7][186] = 1;
   assign ecchmatrix[8][186] = 1;
   assign ecchmatrix[0][187] = 0;
   assign ecchmatrix[1][187] = 1;
   assign ecchmatrix[2][187] = 0;
   assign ecchmatrix[3][187] = 0;
   assign ecchmatrix[4][187] = 1;
   assign ecchmatrix[5][187] = 0;
   assign ecchmatrix[6][187] = 1;
   assign ecchmatrix[7][187] = 1;
   assign ecchmatrix[8][187] = 1;
   assign ecchmatrix[0][188] = 0;
   assign ecchmatrix[1][188] = 1;
   assign ecchmatrix[2][188] = 0;
   assign ecchmatrix[3][188] = 0;
   assign ecchmatrix[4][188] = 0;
   assign ecchmatrix[5][188] = 1;
   assign ecchmatrix[6][188] = 1;
   assign ecchmatrix[7][188] = 1;
   assign ecchmatrix[8][188] = 1;
   assign ecchmatrix[0][189] = 0;
   assign ecchmatrix[1][189] = 0;
   assign ecchmatrix[2][189] = 1;
   assign ecchmatrix[3][189] = 1;
   assign ecchmatrix[4][189] = 1;
   assign ecchmatrix[5][189] = 1;
   assign ecchmatrix[6][189] = 1;
   assign ecchmatrix[7][189] = 0;
   assign ecchmatrix[8][189] = 0;
   assign ecchmatrix[0][190] = 0;
   assign ecchmatrix[1][190] = 0;
   assign ecchmatrix[2][190] = 1;
   assign ecchmatrix[3][190] = 1;
   assign ecchmatrix[4][190] = 1;
   assign ecchmatrix[5][190] = 1;
   assign ecchmatrix[6][190] = 0;
   assign ecchmatrix[7][190] = 1;
   assign ecchmatrix[8][190] = 0;
   assign ecchmatrix[0][191] = 0;
   assign ecchmatrix[1][191] = 0;
   assign ecchmatrix[2][191] = 1;
   assign ecchmatrix[3][191] = 1;
   assign ecchmatrix[4][191] = 1;
   assign ecchmatrix[5][191] = 1;
   assign ecchmatrix[6][191] = 0;
   assign ecchmatrix[7][191] = 0;
   assign ecchmatrix[8][191] = 1;
   assign ecchmatrix[0][192] = 0;
   assign ecchmatrix[1][192] = 0;
   assign ecchmatrix[2][192] = 1;
   assign ecchmatrix[3][192] = 1;
   assign ecchmatrix[4][192] = 1;
   assign ecchmatrix[5][192] = 0;
   assign ecchmatrix[6][192] = 1;
   assign ecchmatrix[7][192] = 1;
   assign ecchmatrix[8][192] = 0;
   assign ecchmatrix[0][193] = 0;
   assign ecchmatrix[1][193] = 0;
   assign ecchmatrix[2][193] = 1;
   assign ecchmatrix[3][193] = 1;
   assign ecchmatrix[4][193] = 1;
   assign ecchmatrix[5][193] = 0;
   assign ecchmatrix[6][193] = 1;
   assign ecchmatrix[7][193] = 0;
   assign ecchmatrix[8][193] = 1;
   assign ecchmatrix[0][194] = 0;
   assign ecchmatrix[1][194] = 0;
   assign ecchmatrix[2][194] = 1;
   assign ecchmatrix[3][194] = 1;
   assign ecchmatrix[4][194] = 1;
   assign ecchmatrix[5][194] = 0;
   assign ecchmatrix[6][194] = 0;
   assign ecchmatrix[7][194] = 1;
   assign ecchmatrix[8][194] = 1;
   assign ecchmatrix[0][195] = 0;
   assign ecchmatrix[1][195] = 0;
   assign ecchmatrix[2][195] = 1;
   assign ecchmatrix[3][195] = 1;
   assign ecchmatrix[4][195] = 0;
   assign ecchmatrix[5][195] = 1;
   assign ecchmatrix[6][195] = 1;
   assign ecchmatrix[7][195] = 1;
   assign ecchmatrix[8][195] = 0;
   assign ecchmatrix[0][196] = 0;
   assign ecchmatrix[1][196] = 0;
   assign ecchmatrix[2][196] = 1;
   assign ecchmatrix[3][196] = 1;
   assign ecchmatrix[4][196] = 0;
   assign ecchmatrix[5][196] = 1;
   assign ecchmatrix[6][196] = 1;
   assign ecchmatrix[7][196] = 0;
   assign ecchmatrix[8][196] = 1;
   assign ecchmatrix[0][197] = 0;
   assign ecchmatrix[1][197] = 0;
   assign ecchmatrix[2][197] = 1;
   assign ecchmatrix[3][197] = 1;
   assign ecchmatrix[4][197] = 0;
   assign ecchmatrix[5][197] = 1;
   assign ecchmatrix[6][197] = 0;
   assign ecchmatrix[7][197] = 1;
   assign ecchmatrix[8][197] = 1;
   assign ecchmatrix[0][198] = 0;
   assign ecchmatrix[1][198] = 0;
   assign ecchmatrix[2][198] = 1;
   assign ecchmatrix[3][198] = 1;
   assign ecchmatrix[4][198] = 0;
   assign ecchmatrix[5][198] = 0;
   assign ecchmatrix[6][198] = 1;
   assign ecchmatrix[7][198] = 1;
   assign ecchmatrix[8][198] = 1;
   assign ecchmatrix[0][199] = 0;
   assign ecchmatrix[1][199] = 0;
   assign ecchmatrix[2][199] = 1;
   assign ecchmatrix[3][199] = 0;
   assign ecchmatrix[4][199] = 1;
   assign ecchmatrix[5][199] = 1;
   assign ecchmatrix[6][199] = 1;
   assign ecchmatrix[7][199] = 1;
   assign ecchmatrix[8][199] = 0;
   assign ecchmatrix[0][200] = 0;
   assign ecchmatrix[1][200] = 0;
   assign ecchmatrix[2][200] = 1;
   assign ecchmatrix[3][200] = 0;
   assign ecchmatrix[4][200] = 1;
   assign ecchmatrix[5][200] = 1;
   assign ecchmatrix[6][200] = 1;
   assign ecchmatrix[7][200] = 0;
   assign ecchmatrix[8][200] = 1;
   assign ecchmatrix[0][201] = 0;
   assign ecchmatrix[1][201] = 0;
   assign ecchmatrix[2][201] = 1;
   assign ecchmatrix[3][201] = 0;
   assign ecchmatrix[4][201] = 1;
   assign ecchmatrix[5][201] = 1;
   assign ecchmatrix[6][201] = 0;
   assign ecchmatrix[7][201] = 1;
   assign ecchmatrix[8][201] = 1;
   assign ecchmatrix[0][202] = 0;
   assign ecchmatrix[1][202] = 0;
   assign ecchmatrix[2][202] = 1;
   assign ecchmatrix[3][202] = 0;
   assign ecchmatrix[4][202] = 1;
   assign ecchmatrix[5][202] = 0;
   assign ecchmatrix[6][202] = 1;
   assign ecchmatrix[7][202] = 1;
   assign ecchmatrix[8][202] = 1;
   assign ecchmatrix[0][203] = 0;
   assign ecchmatrix[1][203] = 0;
   assign ecchmatrix[2][203] = 1;
   assign ecchmatrix[3][203] = 0;
   assign ecchmatrix[4][203] = 0;
   assign ecchmatrix[5][203] = 1;
   assign ecchmatrix[6][203] = 1;
   assign ecchmatrix[7][203] = 1;
   assign ecchmatrix[8][203] = 1;
   assign ecchmatrix[0][204] = 0;
   assign ecchmatrix[1][204] = 0;
   assign ecchmatrix[2][204] = 0;
   assign ecchmatrix[3][204] = 1;
   assign ecchmatrix[4][204] = 1;
   assign ecchmatrix[5][204] = 1;
   assign ecchmatrix[6][204] = 1;
   assign ecchmatrix[7][204] = 1;
   assign ecchmatrix[8][204] = 0;
   assign ecchmatrix[0][205] = 0;
   assign ecchmatrix[1][205] = 0;
   assign ecchmatrix[2][205] = 0;
   assign ecchmatrix[3][205] = 1;
   assign ecchmatrix[4][205] = 1;
   assign ecchmatrix[5][205] = 1;
   assign ecchmatrix[6][205] = 1;
   assign ecchmatrix[7][205] = 0;
   assign ecchmatrix[8][205] = 1;
   assign ecchmatrix[0][206] = 0;
   assign ecchmatrix[1][206] = 0;
   assign ecchmatrix[2][206] = 0;
   assign ecchmatrix[3][206] = 1;
   assign ecchmatrix[4][206] = 1;
   assign ecchmatrix[5][206] = 1;
   assign ecchmatrix[6][206] = 0;
   assign ecchmatrix[7][206] = 1;
   assign ecchmatrix[8][206] = 1;
   assign ecchmatrix[0][207] = 0;
   assign ecchmatrix[1][207] = 0;
   assign ecchmatrix[2][207] = 0;
   assign ecchmatrix[3][207] = 1;
   assign ecchmatrix[4][207] = 1;
   assign ecchmatrix[5][207] = 0;
   assign ecchmatrix[6][207] = 1;
   assign ecchmatrix[7][207] = 1;
   assign ecchmatrix[8][207] = 1;
   assign ecchmatrix[0][208] = 0;
   assign ecchmatrix[1][208] = 0;
   assign ecchmatrix[2][208] = 0;
   assign ecchmatrix[3][208] = 1;
   assign ecchmatrix[4][208] = 0;
   assign ecchmatrix[5][208] = 1;
   assign ecchmatrix[6][208] = 1;
   assign ecchmatrix[7][208] = 1;
   assign ecchmatrix[8][208] = 1;
   assign ecchmatrix[0][209] = 0;
   assign ecchmatrix[1][209] = 0;
   assign ecchmatrix[2][209] = 0;
   assign ecchmatrix[3][209] = 0;
   assign ecchmatrix[4][209] = 1;
   assign ecchmatrix[5][209] = 1;
   assign ecchmatrix[6][209] = 1;
   assign ecchmatrix[7][209] = 1;
   assign ecchmatrix[8][209] = 1;
   assign ecchmatrix[0][210] = 1;
   assign ecchmatrix[1][210] = 1;
   assign ecchmatrix[2][210] = 1;
   assign ecchmatrix[3][210] = 1;
   assign ecchmatrix[4][210] = 1;
   assign ecchmatrix[5][210] = 1;
   assign ecchmatrix[6][210] = 1;
   assign ecchmatrix[7][210] = 0;
   assign ecchmatrix[8][210] = 0;
   assign ecchmatrix[0][211] = 1;
   assign ecchmatrix[1][211] = 1;
   assign ecchmatrix[2][211] = 1;
   assign ecchmatrix[3][211] = 1;
   assign ecchmatrix[4][211] = 1;
   assign ecchmatrix[5][211] = 1;
   assign ecchmatrix[6][211] = 0;
   assign ecchmatrix[7][211] = 1;
   assign ecchmatrix[8][211] = 0;
   assign ecchmatrix[0][212] = 1;
   assign ecchmatrix[1][212] = 1;
   assign ecchmatrix[2][212] = 1;
   assign ecchmatrix[3][212] = 1;
   assign ecchmatrix[4][212] = 1;
   assign ecchmatrix[5][212] = 1;
   assign ecchmatrix[6][212] = 0;
   assign ecchmatrix[7][212] = 0;
   assign ecchmatrix[8][212] = 1;
   assign ecchmatrix[0][213] = 1;
   assign ecchmatrix[1][213] = 1;
   assign ecchmatrix[2][213] = 1;
   assign ecchmatrix[3][213] = 1;
   assign ecchmatrix[4][213] = 1;
   assign ecchmatrix[5][213] = 0;
   assign ecchmatrix[6][213] = 1;
   assign ecchmatrix[7][213] = 1;
   assign ecchmatrix[8][213] = 0;
   assign ecchmatrix[0][214] = 1;
   assign ecchmatrix[1][214] = 1;
   assign ecchmatrix[2][214] = 1;
   assign ecchmatrix[3][214] = 1;
   assign ecchmatrix[4][214] = 1;
   assign ecchmatrix[5][214] = 0;
   assign ecchmatrix[6][214] = 1;
   assign ecchmatrix[7][214] = 0;
   assign ecchmatrix[8][214] = 1;
   assign ecchmatrix[0][215] = 1;
   assign ecchmatrix[1][215] = 1;
   assign ecchmatrix[2][215] = 1;
   assign ecchmatrix[3][215] = 1;
   assign ecchmatrix[4][215] = 1;
   assign ecchmatrix[5][215] = 0;
   assign ecchmatrix[6][215] = 0;
   assign ecchmatrix[7][215] = 1;
   assign ecchmatrix[8][215] = 1;
   assign ecchmatrix[0][216] = 1;
   assign ecchmatrix[1][216] = 1;
   assign ecchmatrix[2][216] = 1;
   assign ecchmatrix[3][216] = 1;
   assign ecchmatrix[4][216] = 0;
   assign ecchmatrix[5][216] = 1;
   assign ecchmatrix[6][216] = 1;
   assign ecchmatrix[7][216] = 1;
   assign ecchmatrix[8][216] = 0;
   assign ecchmatrix[0][217] = 1;
   assign ecchmatrix[1][217] = 1;
   assign ecchmatrix[2][217] = 1;
   assign ecchmatrix[3][217] = 1;
   assign ecchmatrix[4][217] = 0;
   assign ecchmatrix[5][217] = 1;
   assign ecchmatrix[6][217] = 1;
   assign ecchmatrix[7][217] = 0;
   assign ecchmatrix[8][217] = 1;
   assign ecchmatrix[0][218] = 1;
   assign ecchmatrix[1][218] = 1;
   assign ecchmatrix[2][218] = 1;
   assign ecchmatrix[3][218] = 1;
   assign ecchmatrix[4][218] = 0;
   assign ecchmatrix[5][218] = 1;
   assign ecchmatrix[6][218] = 0;
   assign ecchmatrix[7][218] = 1;
   assign ecchmatrix[8][218] = 1;
   assign ecchmatrix[0][219] = 1;
   assign ecchmatrix[1][219] = 1;
   assign ecchmatrix[2][219] = 1;
   assign ecchmatrix[3][219] = 1;
   assign ecchmatrix[4][219] = 0;
   assign ecchmatrix[5][219] = 0;
   assign ecchmatrix[6][219] = 1;
   assign ecchmatrix[7][219] = 1;
   assign ecchmatrix[8][219] = 1;
   assign ecchmatrix[0][220] = 1;
   assign ecchmatrix[1][220] = 1;
   assign ecchmatrix[2][220] = 1;
   assign ecchmatrix[3][220] = 0;
   assign ecchmatrix[4][220] = 1;
   assign ecchmatrix[5][220] = 1;
   assign ecchmatrix[6][220] = 1;
   assign ecchmatrix[7][220] = 1;
   assign ecchmatrix[8][220] = 0;
   assign ecchmatrix[0][221] = 1;
   assign ecchmatrix[1][221] = 1;
   assign ecchmatrix[2][221] = 1;
   assign ecchmatrix[3][221] = 0;
   assign ecchmatrix[4][221] = 1;
   assign ecchmatrix[5][221] = 1;
   assign ecchmatrix[6][221] = 1;
   assign ecchmatrix[7][221] = 0;
   assign ecchmatrix[8][221] = 1;
   assign ecchmatrix[0][222] = 1;
   assign ecchmatrix[1][222] = 1;
   assign ecchmatrix[2][222] = 1;
   assign ecchmatrix[3][222] = 0;
   assign ecchmatrix[4][222] = 1;
   assign ecchmatrix[5][222] = 1;
   assign ecchmatrix[6][222] = 0;
   assign ecchmatrix[7][222] = 1;
   assign ecchmatrix[8][222] = 1;
   assign ecchmatrix[0][223] = 1;
   assign ecchmatrix[1][223] = 1;
   assign ecchmatrix[2][223] = 1;
   assign ecchmatrix[3][223] = 0;
   assign ecchmatrix[4][223] = 1;
   assign ecchmatrix[5][223] = 0;
   assign ecchmatrix[6][223] = 1;
   assign ecchmatrix[7][223] = 1;
   assign ecchmatrix[8][223] = 1;
   assign ecchmatrix[0][224] = 1;
   assign ecchmatrix[1][224] = 1;
   assign ecchmatrix[2][224] = 1;
   assign ecchmatrix[3][224] = 0;
   assign ecchmatrix[4][224] = 0;
   assign ecchmatrix[5][224] = 1;
   assign ecchmatrix[6][224] = 1;
   assign ecchmatrix[7][224] = 1;
   assign ecchmatrix[8][224] = 1;
   assign ecchmatrix[0][225] = 1;
   assign ecchmatrix[1][225] = 1;
   assign ecchmatrix[2][225] = 0;
   assign ecchmatrix[3][225] = 1;
   assign ecchmatrix[4][225] = 1;
   assign ecchmatrix[5][225] = 1;
   assign ecchmatrix[6][225] = 1;
   assign ecchmatrix[7][225] = 1;
   assign ecchmatrix[8][225] = 0;
   assign ecchmatrix[0][226] = 1;
   assign ecchmatrix[1][226] = 1;
   assign ecchmatrix[2][226] = 0;
   assign ecchmatrix[3][226] = 1;
   assign ecchmatrix[4][226] = 1;
   assign ecchmatrix[5][226] = 1;
   assign ecchmatrix[6][226] = 1;
   assign ecchmatrix[7][226] = 0;
   assign ecchmatrix[8][226] = 1;
   assign ecchmatrix[0][227] = 1;
   assign ecchmatrix[1][227] = 1;
   assign ecchmatrix[2][227] = 0;
   assign ecchmatrix[3][227] = 1;
   assign ecchmatrix[4][227] = 1;
   assign ecchmatrix[5][227] = 1;
   assign ecchmatrix[6][227] = 0;
   assign ecchmatrix[7][227] = 1;
   assign ecchmatrix[8][227] = 1;
   assign ecchmatrix[0][228] = 1;
   assign ecchmatrix[1][228] = 1;
   assign ecchmatrix[2][228] = 0;
   assign ecchmatrix[3][228] = 1;
   assign ecchmatrix[4][228] = 1;
   assign ecchmatrix[5][228] = 0;
   assign ecchmatrix[6][228] = 1;
   assign ecchmatrix[7][228] = 1;
   assign ecchmatrix[8][228] = 1;
   assign ecchmatrix[0][229] = 1;
   assign ecchmatrix[1][229] = 1;
   assign ecchmatrix[2][229] = 0;
   assign ecchmatrix[3][229] = 1;
   assign ecchmatrix[4][229] = 0;
   assign ecchmatrix[5][229] = 1;
   assign ecchmatrix[6][229] = 1;
   assign ecchmatrix[7][229] = 1;
   assign ecchmatrix[8][229] = 1;
   assign ecchmatrix[0][230] = 1;
   assign ecchmatrix[1][230] = 1;
   assign ecchmatrix[2][230] = 0;
   assign ecchmatrix[3][230] = 0;
   assign ecchmatrix[4][230] = 1;
   assign ecchmatrix[5][230] = 1;
   assign ecchmatrix[6][230] = 1;
   assign ecchmatrix[7][230] = 1;
   assign ecchmatrix[8][230] = 1;
   assign ecchmatrix[0][231] = 1;
   assign ecchmatrix[1][231] = 0;
   assign ecchmatrix[2][231] = 1;
   assign ecchmatrix[3][231] = 1;
   assign ecchmatrix[4][231] = 1;
   assign ecchmatrix[5][231] = 1;
   assign ecchmatrix[6][231] = 1;
   assign ecchmatrix[7][231] = 1;
   assign ecchmatrix[8][231] = 0;
   assign ecchmatrix[0][232] = 1;
   assign ecchmatrix[1][232] = 0;
   assign ecchmatrix[2][232] = 1;
   assign ecchmatrix[3][232] = 1;
   assign ecchmatrix[4][232] = 1;
   assign ecchmatrix[5][232] = 1;
   assign ecchmatrix[6][232] = 1;
   assign ecchmatrix[7][232] = 0;
   assign ecchmatrix[8][232] = 1;
   assign ecchmatrix[0][233] = 1;
   assign ecchmatrix[1][233] = 0;
   assign ecchmatrix[2][233] = 1;
   assign ecchmatrix[3][233] = 1;
   assign ecchmatrix[4][233] = 1;
   assign ecchmatrix[5][233] = 1;
   assign ecchmatrix[6][233] = 0;
   assign ecchmatrix[7][233] = 1;
   assign ecchmatrix[8][233] = 1;
   assign ecchmatrix[0][234] = 1;
   assign ecchmatrix[1][234] = 0;
   assign ecchmatrix[2][234] = 1;
   assign ecchmatrix[3][234] = 1;
   assign ecchmatrix[4][234] = 1;
   assign ecchmatrix[5][234] = 0;
   assign ecchmatrix[6][234] = 1;
   assign ecchmatrix[7][234] = 1;
   assign ecchmatrix[8][234] = 1;
   assign ecchmatrix[0][235] = 1;
   assign ecchmatrix[1][235] = 0;
   assign ecchmatrix[2][235] = 1;
   assign ecchmatrix[3][235] = 1;
   assign ecchmatrix[4][235] = 0;
   assign ecchmatrix[5][235] = 1;
   assign ecchmatrix[6][235] = 1;
   assign ecchmatrix[7][235] = 1;
   assign ecchmatrix[8][235] = 1;
   assign ecchmatrix[0][236] = 1;
   assign ecchmatrix[1][236] = 0;
   assign ecchmatrix[2][236] = 1;
   assign ecchmatrix[3][236] = 0;
   assign ecchmatrix[4][236] = 1;
   assign ecchmatrix[5][236] = 1;
   assign ecchmatrix[6][236] = 1;
   assign ecchmatrix[7][236] = 1;
   assign ecchmatrix[8][236] = 1;
   assign ecchmatrix[0][237] = 1;
   assign ecchmatrix[1][237] = 0;
   assign ecchmatrix[2][237] = 0;
   assign ecchmatrix[3][237] = 1;
   assign ecchmatrix[4][237] = 1;
   assign ecchmatrix[5][237] = 1;
   assign ecchmatrix[6][237] = 1;
   assign ecchmatrix[7][237] = 1;
   assign ecchmatrix[8][237] = 1;
   assign ecchmatrix[0][238] = 0;
   assign ecchmatrix[1][238] = 1;
   assign ecchmatrix[2][238] = 1;
   assign ecchmatrix[3][238] = 1;
   assign ecchmatrix[4][238] = 1;
   assign ecchmatrix[5][238] = 1;
   assign ecchmatrix[6][238] = 1;
   assign ecchmatrix[7][238] = 1;
   assign ecchmatrix[8][238] = 0;
   assign ecchmatrix[0][239] = 0;
   assign ecchmatrix[1][239] = 1;
   assign ecchmatrix[2][239] = 1;
   assign ecchmatrix[3][239] = 1;
   assign ecchmatrix[4][239] = 1;
   assign ecchmatrix[5][239] = 1;
   assign ecchmatrix[6][239] = 1;
   assign ecchmatrix[7][239] = 0;
   assign ecchmatrix[8][239] = 1;
   assign ecchmatrix[0][240] = 0;
   assign ecchmatrix[1][240] = 1;
   assign ecchmatrix[2][240] = 1;
   assign ecchmatrix[3][240] = 1;
   assign ecchmatrix[4][240] = 1;
   assign ecchmatrix[5][240] = 1;
   assign ecchmatrix[6][240] = 0;
   assign ecchmatrix[7][240] = 1;
   assign ecchmatrix[8][240] = 1;
   assign ecchmatrix[0][241] = 0;
   assign ecchmatrix[1][241] = 1;
   assign ecchmatrix[2][241] = 1;
   assign ecchmatrix[3][241] = 1;
   assign ecchmatrix[4][241] = 1;
   assign ecchmatrix[5][241] = 0;
   assign ecchmatrix[6][241] = 1;
   assign ecchmatrix[7][241] = 1;
   assign ecchmatrix[8][241] = 1;
   assign ecchmatrix[0][242] = 0;
   assign ecchmatrix[1][242] = 1;
   assign ecchmatrix[2][242] = 1;
   assign ecchmatrix[3][242] = 1;
   assign ecchmatrix[4][242] = 0;
   assign ecchmatrix[5][242] = 1;
   assign ecchmatrix[6][242] = 1;
   assign ecchmatrix[7][242] = 1;
   assign ecchmatrix[8][242] = 1;
   assign ecchmatrix[0][243] = 0;
   assign ecchmatrix[1][243] = 1;
   assign ecchmatrix[2][243] = 1;
   assign ecchmatrix[3][243] = 0;
   assign ecchmatrix[4][243] = 1;
   assign ecchmatrix[5][243] = 1;
   assign ecchmatrix[6][243] = 1;
   assign ecchmatrix[7][243] = 1;
   assign ecchmatrix[8][243] = 1;
   assign ecchmatrix[0][244] = 0;
   assign ecchmatrix[1][244] = 1;
   assign ecchmatrix[2][244] = 0;
   assign ecchmatrix[3][244] = 1;
   assign ecchmatrix[4][244] = 1;
   assign ecchmatrix[5][244] = 1;
   assign ecchmatrix[6][244] = 1;
   assign ecchmatrix[7][244] = 1;
   assign ecchmatrix[8][244] = 1;
   assign ecchmatrix[0][245] = 0;
   assign ecchmatrix[1][245] = 0;
   assign ecchmatrix[2][245] = 1;
   assign ecchmatrix[3][245] = 1;
   assign ecchmatrix[4][245] = 1;
   assign ecchmatrix[5][245] = 1;
   assign ecchmatrix[6][245] = 1;
   assign ecchmatrix[7][245] = 1;
   assign ecchmatrix[8][245] = 1;
   assign ecchmatrix[0][246] = 1;
   assign ecchmatrix[1][246] = 1;
   assign ecchmatrix[2][246] = 1;
   assign ecchmatrix[3][246] = 1;
   assign ecchmatrix[4][246] = 1;
   assign ecchmatrix[5][246] = 1;
   assign ecchmatrix[6][246] = 1;
   assign ecchmatrix[7][246] = 1;
   assign ecchmatrix[8][246] = 1;
endmodule

module ecc_calc_502 (din, eccout);

  localparam ECCDWIDTH = 502;
  localparam ECCWIDTH  = 10;
  
  input [ECCDWIDTH-1:0]            din;  
  output [ECCWIDTH-1:0]            eccout;

  wire [ECCDWIDTH-1:0]   ecchmatrix [0:ECCWIDTH-1];

 assign eccout[9] = ^(ecchmatrix[9]&din);
 assign eccout[8] = ^(ecchmatrix[8]&din);
 assign eccout[7] = ^(ecchmatrix[7]&din);
 assign eccout[6] = ^(ecchmatrix[6]&din);
 assign eccout[5] = ^(ecchmatrix[5]&din);
 assign eccout[4] = ^(ecchmatrix[4]&din);
 assign eccout[3] = ^(ecchmatrix[3]&din);
 assign eccout[2] = ^(ecchmatrix[2]&din);
 assign eccout[1] = ^(ecchmatrix[1]&din);
 assign eccout[0] = ^(ecchmatrix[0]&din);
// assign ready = 1'b1;

// Generate the H Matrix in Perl

// Initialize the hmatrix array
   assign ecchmatrix[0][0] = 1;
   assign ecchmatrix[1][0] = 1;
   assign ecchmatrix[2][0] = 1;
   assign ecchmatrix[3][0] = 0;
   assign ecchmatrix[4][0] = 0;
   assign ecchmatrix[5][0] = 0;
   assign ecchmatrix[6][0] = 0;
   assign ecchmatrix[7][0] = 0;
   assign ecchmatrix[8][0] = 0;
   assign ecchmatrix[9][0] = 0;
   assign ecchmatrix[0][1] = 1;
   assign ecchmatrix[1][1] = 1;
   assign ecchmatrix[2][1] = 0;
   assign ecchmatrix[3][1] = 1;
   assign ecchmatrix[4][1] = 0;
   assign ecchmatrix[5][1] = 0;
   assign ecchmatrix[6][1] = 0;
   assign ecchmatrix[7][1] = 0;
   assign ecchmatrix[8][1] = 0;
   assign ecchmatrix[9][1] = 0;
   assign ecchmatrix[0][2] = 1;
   assign ecchmatrix[1][2] = 1;
   assign ecchmatrix[2][2] = 0;
   assign ecchmatrix[3][2] = 0;
   assign ecchmatrix[4][2] = 1;
   assign ecchmatrix[5][2] = 0;
   assign ecchmatrix[6][2] = 0;
   assign ecchmatrix[7][2] = 0;
   assign ecchmatrix[8][2] = 0;
   assign ecchmatrix[9][2] = 0;
   assign ecchmatrix[0][3] = 1;
   assign ecchmatrix[1][3] = 1;
   assign ecchmatrix[2][3] = 0;
   assign ecchmatrix[3][3] = 0;
   assign ecchmatrix[4][3] = 0;
   assign ecchmatrix[5][3] = 1;
   assign ecchmatrix[6][3] = 0;
   assign ecchmatrix[7][3] = 0;
   assign ecchmatrix[8][3] = 0;
   assign ecchmatrix[9][3] = 0;
   assign ecchmatrix[0][4] = 1;
   assign ecchmatrix[1][4] = 1;
   assign ecchmatrix[2][4] = 0;
   assign ecchmatrix[3][4] = 0;
   assign ecchmatrix[4][4] = 0;
   assign ecchmatrix[5][4] = 0;
   assign ecchmatrix[6][4] = 1;
   assign ecchmatrix[7][4] = 0;
   assign ecchmatrix[8][4] = 0;
   assign ecchmatrix[9][4] = 0;
   assign ecchmatrix[0][5] = 1;
   assign ecchmatrix[1][5] = 1;
   assign ecchmatrix[2][5] = 0;
   assign ecchmatrix[3][5] = 0;
   assign ecchmatrix[4][5] = 0;
   assign ecchmatrix[5][5] = 0;
   assign ecchmatrix[6][5] = 0;
   assign ecchmatrix[7][5] = 1;
   assign ecchmatrix[8][5] = 0;
   assign ecchmatrix[9][5] = 0;
   assign ecchmatrix[0][6] = 1;
   assign ecchmatrix[1][6] = 1;
   assign ecchmatrix[2][6] = 0;
   assign ecchmatrix[3][6] = 0;
   assign ecchmatrix[4][6] = 0;
   assign ecchmatrix[5][6] = 0;
   assign ecchmatrix[6][6] = 0;
   assign ecchmatrix[7][6] = 0;
   assign ecchmatrix[8][6] = 1;
   assign ecchmatrix[9][6] = 0;
   assign ecchmatrix[0][7] = 1;
   assign ecchmatrix[1][7] = 1;
   assign ecchmatrix[2][7] = 0;
   assign ecchmatrix[3][7] = 0;
   assign ecchmatrix[4][7] = 0;
   assign ecchmatrix[5][7] = 0;
   assign ecchmatrix[6][7] = 0;
   assign ecchmatrix[7][7] = 0;
   assign ecchmatrix[8][7] = 0;
   assign ecchmatrix[9][7] = 1;
   assign ecchmatrix[0][8] = 1;
   assign ecchmatrix[1][8] = 0;
   assign ecchmatrix[2][8] = 1;
   assign ecchmatrix[3][8] = 1;
   assign ecchmatrix[4][8] = 0;
   assign ecchmatrix[5][8] = 0;
   assign ecchmatrix[6][8] = 0;
   assign ecchmatrix[7][8] = 0;
   assign ecchmatrix[8][8] = 0;
   assign ecchmatrix[9][8] = 0;
   assign ecchmatrix[0][9] = 1;
   assign ecchmatrix[1][9] = 0;
   assign ecchmatrix[2][9] = 1;
   assign ecchmatrix[3][9] = 0;
   assign ecchmatrix[4][9] = 1;
   assign ecchmatrix[5][9] = 0;
   assign ecchmatrix[6][9] = 0;
   assign ecchmatrix[7][9] = 0;
   assign ecchmatrix[8][9] = 0;
   assign ecchmatrix[9][9] = 0;
   assign ecchmatrix[0][10] = 1;
   assign ecchmatrix[1][10] = 0;
   assign ecchmatrix[2][10] = 1;
   assign ecchmatrix[3][10] = 0;
   assign ecchmatrix[4][10] = 0;
   assign ecchmatrix[5][10] = 1;
   assign ecchmatrix[6][10] = 0;
   assign ecchmatrix[7][10] = 0;
   assign ecchmatrix[8][10] = 0;
   assign ecchmatrix[9][10] = 0;
   assign ecchmatrix[0][11] = 1;
   assign ecchmatrix[1][11] = 0;
   assign ecchmatrix[2][11] = 1;
   assign ecchmatrix[3][11] = 0;
   assign ecchmatrix[4][11] = 0;
   assign ecchmatrix[5][11] = 0;
   assign ecchmatrix[6][11] = 1;
   assign ecchmatrix[7][11] = 0;
   assign ecchmatrix[8][11] = 0;
   assign ecchmatrix[9][11] = 0;
   assign ecchmatrix[0][12] = 1;
   assign ecchmatrix[1][12] = 0;
   assign ecchmatrix[2][12] = 1;
   assign ecchmatrix[3][12] = 0;
   assign ecchmatrix[4][12] = 0;
   assign ecchmatrix[5][12] = 0;
   assign ecchmatrix[6][12] = 0;
   assign ecchmatrix[7][12] = 1;
   assign ecchmatrix[8][12] = 0;
   assign ecchmatrix[9][12] = 0;
   assign ecchmatrix[0][13] = 1;
   assign ecchmatrix[1][13] = 0;
   assign ecchmatrix[2][13] = 1;
   assign ecchmatrix[3][13] = 0;
   assign ecchmatrix[4][13] = 0;
   assign ecchmatrix[5][13] = 0;
   assign ecchmatrix[6][13] = 0;
   assign ecchmatrix[7][13] = 0;
   assign ecchmatrix[8][13] = 1;
   assign ecchmatrix[9][13] = 0;
   assign ecchmatrix[0][14] = 1;
   assign ecchmatrix[1][14] = 0;
   assign ecchmatrix[2][14] = 1;
   assign ecchmatrix[3][14] = 0;
   assign ecchmatrix[4][14] = 0;
   assign ecchmatrix[5][14] = 0;
   assign ecchmatrix[6][14] = 0;
   assign ecchmatrix[7][14] = 0;
   assign ecchmatrix[8][14] = 0;
   assign ecchmatrix[9][14] = 1;
   assign ecchmatrix[0][15] = 1;
   assign ecchmatrix[1][15] = 0;
   assign ecchmatrix[2][15] = 0;
   assign ecchmatrix[3][15] = 1;
   assign ecchmatrix[4][15] = 1;
   assign ecchmatrix[5][15] = 0;
   assign ecchmatrix[6][15] = 0;
   assign ecchmatrix[7][15] = 0;
   assign ecchmatrix[8][15] = 0;
   assign ecchmatrix[9][15] = 0;
   assign ecchmatrix[0][16] = 1;
   assign ecchmatrix[1][16] = 0;
   assign ecchmatrix[2][16] = 0;
   assign ecchmatrix[3][16] = 1;
   assign ecchmatrix[4][16] = 0;
   assign ecchmatrix[5][16] = 1;
   assign ecchmatrix[6][16] = 0;
   assign ecchmatrix[7][16] = 0;
   assign ecchmatrix[8][16] = 0;
   assign ecchmatrix[9][16] = 0;
   assign ecchmatrix[0][17] = 1;
   assign ecchmatrix[1][17] = 0;
   assign ecchmatrix[2][17] = 0;
   assign ecchmatrix[3][17] = 1;
   assign ecchmatrix[4][17] = 0;
   assign ecchmatrix[5][17] = 0;
   assign ecchmatrix[6][17] = 1;
   assign ecchmatrix[7][17] = 0;
   assign ecchmatrix[8][17] = 0;
   assign ecchmatrix[9][17] = 0;
   assign ecchmatrix[0][18] = 1;
   assign ecchmatrix[1][18] = 0;
   assign ecchmatrix[2][18] = 0;
   assign ecchmatrix[3][18] = 1;
   assign ecchmatrix[4][18] = 0;
   assign ecchmatrix[5][18] = 0;
   assign ecchmatrix[6][18] = 0;
   assign ecchmatrix[7][18] = 1;
   assign ecchmatrix[8][18] = 0;
   assign ecchmatrix[9][18] = 0;
   assign ecchmatrix[0][19] = 1;
   assign ecchmatrix[1][19] = 0;
   assign ecchmatrix[2][19] = 0;
   assign ecchmatrix[3][19] = 1;
   assign ecchmatrix[4][19] = 0;
   assign ecchmatrix[5][19] = 0;
   assign ecchmatrix[6][19] = 0;
   assign ecchmatrix[7][19] = 0;
   assign ecchmatrix[8][19] = 1;
   assign ecchmatrix[9][19] = 0;
   assign ecchmatrix[0][20] = 1;
   assign ecchmatrix[1][20] = 0;
   assign ecchmatrix[2][20] = 0;
   assign ecchmatrix[3][20] = 1;
   assign ecchmatrix[4][20] = 0;
   assign ecchmatrix[5][20] = 0;
   assign ecchmatrix[6][20] = 0;
   assign ecchmatrix[7][20] = 0;
   assign ecchmatrix[8][20] = 0;
   assign ecchmatrix[9][20] = 1;
   assign ecchmatrix[0][21] = 1;
   assign ecchmatrix[1][21] = 0;
   assign ecchmatrix[2][21] = 0;
   assign ecchmatrix[3][21] = 0;
   assign ecchmatrix[4][21] = 1;
   assign ecchmatrix[5][21] = 1;
   assign ecchmatrix[6][21] = 0;
   assign ecchmatrix[7][21] = 0;
   assign ecchmatrix[8][21] = 0;
   assign ecchmatrix[9][21] = 0;
   assign ecchmatrix[0][22] = 1;
   assign ecchmatrix[1][22] = 0;
   assign ecchmatrix[2][22] = 0;
   assign ecchmatrix[3][22] = 0;
   assign ecchmatrix[4][22] = 1;
   assign ecchmatrix[5][22] = 0;
   assign ecchmatrix[6][22] = 1;
   assign ecchmatrix[7][22] = 0;
   assign ecchmatrix[8][22] = 0;
   assign ecchmatrix[9][22] = 0;
   assign ecchmatrix[0][23] = 1;
   assign ecchmatrix[1][23] = 0;
   assign ecchmatrix[2][23] = 0;
   assign ecchmatrix[3][23] = 0;
   assign ecchmatrix[4][23] = 1;
   assign ecchmatrix[5][23] = 0;
   assign ecchmatrix[6][23] = 0;
   assign ecchmatrix[7][23] = 1;
   assign ecchmatrix[8][23] = 0;
   assign ecchmatrix[9][23] = 0;
   assign ecchmatrix[0][24] = 1;
   assign ecchmatrix[1][24] = 0;
   assign ecchmatrix[2][24] = 0;
   assign ecchmatrix[3][24] = 0;
   assign ecchmatrix[4][24] = 1;
   assign ecchmatrix[5][24] = 0;
   assign ecchmatrix[6][24] = 0;
   assign ecchmatrix[7][24] = 0;
   assign ecchmatrix[8][24] = 1;
   assign ecchmatrix[9][24] = 0;
   assign ecchmatrix[0][25] = 1;
   assign ecchmatrix[1][25] = 0;
   assign ecchmatrix[2][25] = 0;
   assign ecchmatrix[3][25] = 0;
   assign ecchmatrix[4][25] = 1;
   assign ecchmatrix[5][25] = 0;
   assign ecchmatrix[6][25] = 0;
   assign ecchmatrix[7][25] = 0;
   assign ecchmatrix[8][25] = 0;
   assign ecchmatrix[9][25] = 1;
   assign ecchmatrix[0][26] = 1;
   assign ecchmatrix[1][26] = 0;
   assign ecchmatrix[2][26] = 0;
   assign ecchmatrix[3][26] = 0;
   assign ecchmatrix[4][26] = 0;
   assign ecchmatrix[5][26] = 1;
   assign ecchmatrix[6][26] = 1;
   assign ecchmatrix[7][26] = 0;
   assign ecchmatrix[8][26] = 0;
   assign ecchmatrix[9][26] = 0;
   assign ecchmatrix[0][27] = 1;
   assign ecchmatrix[1][27] = 0;
   assign ecchmatrix[2][27] = 0;
   assign ecchmatrix[3][27] = 0;
   assign ecchmatrix[4][27] = 0;
   assign ecchmatrix[5][27] = 1;
   assign ecchmatrix[6][27] = 0;
   assign ecchmatrix[7][27] = 1;
   assign ecchmatrix[8][27] = 0;
   assign ecchmatrix[9][27] = 0;
   assign ecchmatrix[0][28] = 1;
   assign ecchmatrix[1][28] = 0;
   assign ecchmatrix[2][28] = 0;
   assign ecchmatrix[3][28] = 0;
   assign ecchmatrix[4][28] = 0;
   assign ecchmatrix[5][28] = 1;
   assign ecchmatrix[6][28] = 0;
   assign ecchmatrix[7][28] = 0;
   assign ecchmatrix[8][28] = 1;
   assign ecchmatrix[9][28] = 0;
   assign ecchmatrix[0][29] = 1;
   assign ecchmatrix[1][29] = 0;
   assign ecchmatrix[2][29] = 0;
   assign ecchmatrix[3][29] = 0;
   assign ecchmatrix[4][29] = 0;
   assign ecchmatrix[5][29] = 1;
   assign ecchmatrix[6][29] = 0;
   assign ecchmatrix[7][29] = 0;
   assign ecchmatrix[8][29] = 0;
   assign ecchmatrix[9][29] = 1;
   assign ecchmatrix[0][30] = 1;
   assign ecchmatrix[1][30] = 0;
   assign ecchmatrix[2][30] = 0;
   assign ecchmatrix[3][30] = 0;
   assign ecchmatrix[4][30] = 0;
   assign ecchmatrix[5][30] = 0;
   assign ecchmatrix[6][30] = 1;
   assign ecchmatrix[7][30] = 1;
   assign ecchmatrix[8][30] = 0;
   assign ecchmatrix[9][30] = 0;
   assign ecchmatrix[0][31] = 1;
   assign ecchmatrix[1][31] = 0;
   assign ecchmatrix[2][31] = 0;
   assign ecchmatrix[3][31] = 0;
   assign ecchmatrix[4][31] = 0;
   assign ecchmatrix[5][31] = 0;
   assign ecchmatrix[6][31] = 1;
   assign ecchmatrix[7][31] = 0;
   assign ecchmatrix[8][31] = 1;
   assign ecchmatrix[9][31] = 0;
   assign ecchmatrix[0][32] = 1;
   assign ecchmatrix[1][32] = 0;
   assign ecchmatrix[2][32] = 0;
   assign ecchmatrix[3][32] = 0;
   assign ecchmatrix[4][32] = 0;
   assign ecchmatrix[5][32] = 0;
   assign ecchmatrix[6][32] = 1;
   assign ecchmatrix[7][32] = 0;
   assign ecchmatrix[8][32] = 0;
   assign ecchmatrix[9][32] = 1;
   assign ecchmatrix[0][33] = 1;
   assign ecchmatrix[1][33] = 0;
   assign ecchmatrix[2][33] = 0;
   assign ecchmatrix[3][33] = 0;
   assign ecchmatrix[4][33] = 0;
   assign ecchmatrix[5][33] = 0;
   assign ecchmatrix[6][33] = 0;
   assign ecchmatrix[7][33] = 1;
   assign ecchmatrix[8][33] = 1;
   assign ecchmatrix[9][33] = 0;
   assign ecchmatrix[0][34] = 1;
   assign ecchmatrix[1][34] = 0;
   assign ecchmatrix[2][34] = 0;
   assign ecchmatrix[3][34] = 0;
   assign ecchmatrix[4][34] = 0;
   assign ecchmatrix[5][34] = 0;
   assign ecchmatrix[6][34] = 0;
   assign ecchmatrix[7][34] = 1;
   assign ecchmatrix[8][34] = 0;
   assign ecchmatrix[9][34] = 1;
   assign ecchmatrix[0][35] = 1;
   assign ecchmatrix[1][35] = 0;
   assign ecchmatrix[2][35] = 0;
   assign ecchmatrix[3][35] = 0;
   assign ecchmatrix[4][35] = 0;
   assign ecchmatrix[5][35] = 0;
   assign ecchmatrix[6][35] = 0;
   assign ecchmatrix[7][35] = 0;
   assign ecchmatrix[8][35] = 1;
   assign ecchmatrix[9][35] = 1;
   assign ecchmatrix[0][36] = 0;
   assign ecchmatrix[1][36] = 1;
   assign ecchmatrix[2][36] = 1;
   assign ecchmatrix[3][36] = 1;
   assign ecchmatrix[4][36] = 0;
   assign ecchmatrix[5][36] = 0;
   assign ecchmatrix[6][36] = 0;
   assign ecchmatrix[7][36] = 0;
   assign ecchmatrix[8][36] = 0;
   assign ecchmatrix[9][36] = 0;
   assign ecchmatrix[0][37] = 0;
   assign ecchmatrix[1][37] = 1;
   assign ecchmatrix[2][37] = 1;
   assign ecchmatrix[3][37] = 0;
   assign ecchmatrix[4][37] = 1;
   assign ecchmatrix[5][37] = 0;
   assign ecchmatrix[6][37] = 0;
   assign ecchmatrix[7][37] = 0;
   assign ecchmatrix[8][37] = 0;
   assign ecchmatrix[9][37] = 0;
   assign ecchmatrix[0][38] = 0;
   assign ecchmatrix[1][38] = 1;
   assign ecchmatrix[2][38] = 1;
   assign ecchmatrix[3][38] = 0;
   assign ecchmatrix[4][38] = 0;
   assign ecchmatrix[5][38] = 1;
   assign ecchmatrix[6][38] = 0;
   assign ecchmatrix[7][38] = 0;
   assign ecchmatrix[8][38] = 0;
   assign ecchmatrix[9][38] = 0;
   assign ecchmatrix[0][39] = 0;
   assign ecchmatrix[1][39] = 1;
   assign ecchmatrix[2][39] = 1;
   assign ecchmatrix[3][39] = 0;
   assign ecchmatrix[4][39] = 0;
   assign ecchmatrix[5][39] = 0;
   assign ecchmatrix[6][39] = 1;
   assign ecchmatrix[7][39] = 0;
   assign ecchmatrix[8][39] = 0;
   assign ecchmatrix[9][39] = 0;
   assign ecchmatrix[0][40] = 0;
   assign ecchmatrix[1][40] = 1;
   assign ecchmatrix[2][40] = 1;
   assign ecchmatrix[3][40] = 0;
   assign ecchmatrix[4][40] = 0;
   assign ecchmatrix[5][40] = 0;
   assign ecchmatrix[6][40] = 0;
   assign ecchmatrix[7][40] = 1;
   assign ecchmatrix[8][40] = 0;
   assign ecchmatrix[9][40] = 0;
   assign ecchmatrix[0][41] = 0;
   assign ecchmatrix[1][41] = 1;
   assign ecchmatrix[2][41] = 1;
   assign ecchmatrix[3][41] = 0;
   assign ecchmatrix[4][41] = 0;
   assign ecchmatrix[5][41] = 0;
   assign ecchmatrix[6][41] = 0;
   assign ecchmatrix[7][41] = 0;
   assign ecchmatrix[8][41] = 1;
   assign ecchmatrix[9][41] = 0;
   assign ecchmatrix[0][42] = 0;
   assign ecchmatrix[1][42] = 1;
   assign ecchmatrix[2][42] = 1;
   assign ecchmatrix[3][42] = 0;
   assign ecchmatrix[4][42] = 0;
   assign ecchmatrix[5][42] = 0;
   assign ecchmatrix[6][42] = 0;
   assign ecchmatrix[7][42] = 0;
   assign ecchmatrix[8][42] = 0;
   assign ecchmatrix[9][42] = 1;
   assign ecchmatrix[0][43] = 0;
   assign ecchmatrix[1][43] = 1;
   assign ecchmatrix[2][43] = 0;
   assign ecchmatrix[3][43] = 1;
   assign ecchmatrix[4][43] = 1;
   assign ecchmatrix[5][43] = 0;
   assign ecchmatrix[6][43] = 0;
   assign ecchmatrix[7][43] = 0;
   assign ecchmatrix[8][43] = 0;
   assign ecchmatrix[9][43] = 0;
   assign ecchmatrix[0][44] = 0;
   assign ecchmatrix[1][44] = 1;
   assign ecchmatrix[2][44] = 0;
   assign ecchmatrix[3][44] = 1;
   assign ecchmatrix[4][44] = 0;
   assign ecchmatrix[5][44] = 1;
   assign ecchmatrix[6][44] = 0;
   assign ecchmatrix[7][44] = 0;
   assign ecchmatrix[8][44] = 0;
   assign ecchmatrix[9][44] = 0;
   assign ecchmatrix[0][45] = 0;
   assign ecchmatrix[1][45] = 1;
   assign ecchmatrix[2][45] = 0;
   assign ecchmatrix[3][45] = 1;
   assign ecchmatrix[4][45] = 0;
   assign ecchmatrix[5][45] = 0;
   assign ecchmatrix[6][45] = 1;
   assign ecchmatrix[7][45] = 0;
   assign ecchmatrix[8][45] = 0;
   assign ecchmatrix[9][45] = 0;
   assign ecchmatrix[0][46] = 0;
   assign ecchmatrix[1][46] = 1;
   assign ecchmatrix[2][46] = 0;
   assign ecchmatrix[3][46] = 1;
   assign ecchmatrix[4][46] = 0;
   assign ecchmatrix[5][46] = 0;
   assign ecchmatrix[6][46] = 0;
   assign ecchmatrix[7][46] = 1;
   assign ecchmatrix[8][46] = 0;
   assign ecchmatrix[9][46] = 0;
   assign ecchmatrix[0][47] = 0;
   assign ecchmatrix[1][47] = 1;
   assign ecchmatrix[2][47] = 0;
   assign ecchmatrix[3][47] = 1;
   assign ecchmatrix[4][47] = 0;
   assign ecchmatrix[5][47] = 0;
   assign ecchmatrix[6][47] = 0;
   assign ecchmatrix[7][47] = 0;
   assign ecchmatrix[8][47] = 1;
   assign ecchmatrix[9][47] = 0;
   assign ecchmatrix[0][48] = 0;
   assign ecchmatrix[1][48] = 1;
   assign ecchmatrix[2][48] = 0;
   assign ecchmatrix[3][48] = 1;
   assign ecchmatrix[4][48] = 0;
   assign ecchmatrix[5][48] = 0;
   assign ecchmatrix[6][48] = 0;
   assign ecchmatrix[7][48] = 0;
   assign ecchmatrix[8][48] = 0;
   assign ecchmatrix[9][48] = 1;
   assign ecchmatrix[0][49] = 0;
   assign ecchmatrix[1][49] = 1;
   assign ecchmatrix[2][49] = 0;
   assign ecchmatrix[3][49] = 0;
   assign ecchmatrix[4][49] = 1;
   assign ecchmatrix[5][49] = 1;
   assign ecchmatrix[6][49] = 0;
   assign ecchmatrix[7][49] = 0;
   assign ecchmatrix[8][49] = 0;
   assign ecchmatrix[9][49] = 0;
   assign ecchmatrix[0][50] = 0;
   assign ecchmatrix[1][50] = 1;
   assign ecchmatrix[2][50] = 0;
   assign ecchmatrix[3][50] = 0;
   assign ecchmatrix[4][50] = 1;
   assign ecchmatrix[5][50] = 0;
   assign ecchmatrix[6][50] = 1;
   assign ecchmatrix[7][50] = 0;
   assign ecchmatrix[8][50] = 0;
   assign ecchmatrix[9][50] = 0;
   assign ecchmatrix[0][51] = 0;
   assign ecchmatrix[1][51] = 1;
   assign ecchmatrix[2][51] = 0;
   assign ecchmatrix[3][51] = 0;
   assign ecchmatrix[4][51] = 1;
   assign ecchmatrix[5][51] = 0;
   assign ecchmatrix[6][51] = 0;
   assign ecchmatrix[7][51] = 1;
   assign ecchmatrix[8][51] = 0;
   assign ecchmatrix[9][51] = 0;
   assign ecchmatrix[0][52] = 0;
   assign ecchmatrix[1][52] = 1;
   assign ecchmatrix[2][52] = 0;
   assign ecchmatrix[3][52] = 0;
   assign ecchmatrix[4][52] = 1;
   assign ecchmatrix[5][52] = 0;
   assign ecchmatrix[6][52] = 0;
   assign ecchmatrix[7][52] = 0;
   assign ecchmatrix[8][52] = 1;
   assign ecchmatrix[9][52] = 0;
   assign ecchmatrix[0][53] = 0;
   assign ecchmatrix[1][53] = 1;
   assign ecchmatrix[2][53] = 0;
   assign ecchmatrix[3][53] = 0;
   assign ecchmatrix[4][53] = 1;
   assign ecchmatrix[5][53] = 0;
   assign ecchmatrix[6][53] = 0;
   assign ecchmatrix[7][53] = 0;
   assign ecchmatrix[8][53] = 0;
   assign ecchmatrix[9][53] = 1;
   assign ecchmatrix[0][54] = 0;
   assign ecchmatrix[1][54] = 1;
   assign ecchmatrix[2][54] = 0;
   assign ecchmatrix[3][54] = 0;
   assign ecchmatrix[4][54] = 0;
   assign ecchmatrix[5][54] = 1;
   assign ecchmatrix[6][54] = 1;
   assign ecchmatrix[7][54] = 0;
   assign ecchmatrix[8][54] = 0;
   assign ecchmatrix[9][54] = 0;
   assign ecchmatrix[0][55] = 0;
   assign ecchmatrix[1][55] = 1;
   assign ecchmatrix[2][55] = 0;
   assign ecchmatrix[3][55] = 0;
   assign ecchmatrix[4][55] = 0;
   assign ecchmatrix[5][55] = 1;
   assign ecchmatrix[6][55] = 0;
   assign ecchmatrix[7][55] = 1;
   assign ecchmatrix[8][55] = 0;
   assign ecchmatrix[9][55] = 0;
   assign ecchmatrix[0][56] = 0;
   assign ecchmatrix[1][56] = 1;
   assign ecchmatrix[2][56] = 0;
   assign ecchmatrix[3][56] = 0;
   assign ecchmatrix[4][56] = 0;
   assign ecchmatrix[5][56] = 1;
   assign ecchmatrix[6][56] = 0;
   assign ecchmatrix[7][56] = 0;
   assign ecchmatrix[8][56] = 1;
   assign ecchmatrix[9][56] = 0;
   assign ecchmatrix[0][57] = 0;
   assign ecchmatrix[1][57] = 1;
   assign ecchmatrix[2][57] = 0;
   assign ecchmatrix[3][57] = 0;
   assign ecchmatrix[4][57] = 0;
   assign ecchmatrix[5][57] = 1;
   assign ecchmatrix[6][57] = 0;
   assign ecchmatrix[7][57] = 0;
   assign ecchmatrix[8][57] = 0;
   assign ecchmatrix[9][57] = 1;
   assign ecchmatrix[0][58] = 0;
   assign ecchmatrix[1][58] = 1;
   assign ecchmatrix[2][58] = 0;
   assign ecchmatrix[3][58] = 0;
   assign ecchmatrix[4][58] = 0;
   assign ecchmatrix[5][58] = 0;
   assign ecchmatrix[6][58] = 1;
   assign ecchmatrix[7][58] = 1;
   assign ecchmatrix[8][58] = 0;
   assign ecchmatrix[9][58] = 0;
   assign ecchmatrix[0][59] = 0;
   assign ecchmatrix[1][59] = 1;
   assign ecchmatrix[2][59] = 0;
   assign ecchmatrix[3][59] = 0;
   assign ecchmatrix[4][59] = 0;
   assign ecchmatrix[5][59] = 0;
   assign ecchmatrix[6][59] = 1;
   assign ecchmatrix[7][59] = 0;
   assign ecchmatrix[8][59] = 1;
   assign ecchmatrix[9][59] = 0;
   assign ecchmatrix[0][60] = 0;
   assign ecchmatrix[1][60] = 1;
   assign ecchmatrix[2][60] = 0;
   assign ecchmatrix[3][60] = 0;
   assign ecchmatrix[4][60] = 0;
   assign ecchmatrix[5][60] = 0;
   assign ecchmatrix[6][60] = 1;
   assign ecchmatrix[7][60] = 0;
   assign ecchmatrix[8][60] = 0;
   assign ecchmatrix[9][60] = 1;
   assign ecchmatrix[0][61] = 0;
   assign ecchmatrix[1][61] = 1;
   assign ecchmatrix[2][61] = 0;
   assign ecchmatrix[3][61] = 0;
   assign ecchmatrix[4][61] = 0;
   assign ecchmatrix[5][61] = 0;
   assign ecchmatrix[6][61] = 0;
   assign ecchmatrix[7][61] = 1;
   assign ecchmatrix[8][61] = 1;
   assign ecchmatrix[9][61] = 0;
   assign ecchmatrix[0][62] = 0;
   assign ecchmatrix[1][62] = 1;
   assign ecchmatrix[2][62] = 0;
   assign ecchmatrix[3][62] = 0;
   assign ecchmatrix[4][62] = 0;
   assign ecchmatrix[5][62] = 0;
   assign ecchmatrix[6][62] = 0;
   assign ecchmatrix[7][62] = 1;
   assign ecchmatrix[8][62] = 0;
   assign ecchmatrix[9][62] = 1;
   assign ecchmatrix[0][63] = 0;
   assign ecchmatrix[1][63] = 1;
   assign ecchmatrix[2][63] = 0;
   assign ecchmatrix[3][63] = 0;
   assign ecchmatrix[4][63] = 0;
   assign ecchmatrix[5][63] = 0;
   assign ecchmatrix[6][63] = 0;
   assign ecchmatrix[7][63] = 0;
   assign ecchmatrix[8][63] = 1;
   assign ecchmatrix[9][63] = 1;
   assign ecchmatrix[0][64] = 0;
   assign ecchmatrix[1][64] = 0;
   assign ecchmatrix[2][64] = 1;
   assign ecchmatrix[3][64] = 1;
   assign ecchmatrix[4][64] = 1;
   assign ecchmatrix[5][64] = 0;
   assign ecchmatrix[6][64] = 0;
   assign ecchmatrix[7][64] = 0;
   assign ecchmatrix[8][64] = 0;
   assign ecchmatrix[9][64] = 0;
   assign ecchmatrix[0][65] = 0;
   assign ecchmatrix[1][65] = 0;
   assign ecchmatrix[2][65] = 1;
   assign ecchmatrix[3][65] = 1;
   assign ecchmatrix[4][65] = 0;
   assign ecchmatrix[5][65] = 1;
   assign ecchmatrix[6][65] = 0;
   assign ecchmatrix[7][65] = 0;
   assign ecchmatrix[8][65] = 0;
   assign ecchmatrix[9][65] = 0;
   assign ecchmatrix[0][66] = 0;
   assign ecchmatrix[1][66] = 0;
   assign ecchmatrix[2][66] = 1;
   assign ecchmatrix[3][66] = 1;
   assign ecchmatrix[4][66] = 0;
   assign ecchmatrix[5][66] = 0;
   assign ecchmatrix[6][66] = 1;
   assign ecchmatrix[7][66] = 0;
   assign ecchmatrix[8][66] = 0;
   assign ecchmatrix[9][66] = 0;
   assign ecchmatrix[0][67] = 0;
   assign ecchmatrix[1][67] = 0;
   assign ecchmatrix[2][67] = 1;
   assign ecchmatrix[3][67] = 1;
   assign ecchmatrix[4][67] = 0;
   assign ecchmatrix[5][67] = 0;
   assign ecchmatrix[6][67] = 0;
   assign ecchmatrix[7][67] = 1;
   assign ecchmatrix[8][67] = 0;
   assign ecchmatrix[9][67] = 0;
   assign ecchmatrix[0][68] = 0;
   assign ecchmatrix[1][68] = 0;
   assign ecchmatrix[2][68] = 1;
   assign ecchmatrix[3][68] = 1;
   assign ecchmatrix[4][68] = 0;
   assign ecchmatrix[5][68] = 0;
   assign ecchmatrix[6][68] = 0;
   assign ecchmatrix[7][68] = 0;
   assign ecchmatrix[8][68] = 1;
   assign ecchmatrix[9][68] = 0;
   assign ecchmatrix[0][69] = 0;
   assign ecchmatrix[1][69] = 0;
   assign ecchmatrix[2][69] = 1;
   assign ecchmatrix[3][69] = 1;
   assign ecchmatrix[4][69] = 0;
   assign ecchmatrix[5][69] = 0;
   assign ecchmatrix[6][69] = 0;
   assign ecchmatrix[7][69] = 0;
   assign ecchmatrix[8][69] = 0;
   assign ecchmatrix[9][69] = 1;
   assign ecchmatrix[0][70] = 0;
   assign ecchmatrix[1][70] = 0;
   assign ecchmatrix[2][70] = 1;
   assign ecchmatrix[3][70] = 0;
   assign ecchmatrix[4][70] = 1;
   assign ecchmatrix[5][70] = 1;
   assign ecchmatrix[6][70] = 0;
   assign ecchmatrix[7][70] = 0;
   assign ecchmatrix[8][70] = 0;
   assign ecchmatrix[9][70] = 0;
   assign ecchmatrix[0][71] = 0;
   assign ecchmatrix[1][71] = 0;
   assign ecchmatrix[2][71] = 1;
   assign ecchmatrix[3][71] = 0;
   assign ecchmatrix[4][71] = 1;
   assign ecchmatrix[5][71] = 0;
   assign ecchmatrix[6][71] = 1;
   assign ecchmatrix[7][71] = 0;
   assign ecchmatrix[8][71] = 0;
   assign ecchmatrix[9][71] = 0;
   assign ecchmatrix[0][72] = 0;
   assign ecchmatrix[1][72] = 0;
   assign ecchmatrix[2][72] = 1;
   assign ecchmatrix[3][72] = 0;
   assign ecchmatrix[4][72] = 1;
   assign ecchmatrix[5][72] = 0;
   assign ecchmatrix[6][72] = 0;
   assign ecchmatrix[7][72] = 1;
   assign ecchmatrix[8][72] = 0;
   assign ecchmatrix[9][72] = 0;
   assign ecchmatrix[0][73] = 0;
   assign ecchmatrix[1][73] = 0;
   assign ecchmatrix[2][73] = 1;
   assign ecchmatrix[3][73] = 0;
   assign ecchmatrix[4][73] = 1;
   assign ecchmatrix[5][73] = 0;
   assign ecchmatrix[6][73] = 0;
   assign ecchmatrix[7][73] = 0;
   assign ecchmatrix[8][73] = 1;
   assign ecchmatrix[9][73] = 0;
   assign ecchmatrix[0][74] = 0;
   assign ecchmatrix[1][74] = 0;
   assign ecchmatrix[2][74] = 1;
   assign ecchmatrix[3][74] = 0;
   assign ecchmatrix[4][74] = 1;
   assign ecchmatrix[5][74] = 0;
   assign ecchmatrix[6][74] = 0;
   assign ecchmatrix[7][74] = 0;
   assign ecchmatrix[8][74] = 0;
   assign ecchmatrix[9][74] = 1;
   assign ecchmatrix[0][75] = 0;
   assign ecchmatrix[1][75] = 0;
   assign ecchmatrix[2][75] = 1;
   assign ecchmatrix[3][75] = 0;
   assign ecchmatrix[4][75] = 0;
   assign ecchmatrix[5][75] = 1;
   assign ecchmatrix[6][75] = 1;
   assign ecchmatrix[7][75] = 0;
   assign ecchmatrix[8][75] = 0;
   assign ecchmatrix[9][75] = 0;
   assign ecchmatrix[0][76] = 0;
   assign ecchmatrix[1][76] = 0;
   assign ecchmatrix[2][76] = 1;
   assign ecchmatrix[3][76] = 0;
   assign ecchmatrix[4][76] = 0;
   assign ecchmatrix[5][76] = 1;
   assign ecchmatrix[6][76] = 0;
   assign ecchmatrix[7][76] = 1;
   assign ecchmatrix[8][76] = 0;
   assign ecchmatrix[9][76] = 0;
   assign ecchmatrix[0][77] = 0;
   assign ecchmatrix[1][77] = 0;
   assign ecchmatrix[2][77] = 1;
   assign ecchmatrix[3][77] = 0;
   assign ecchmatrix[4][77] = 0;
   assign ecchmatrix[5][77] = 1;
   assign ecchmatrix[6][77] = 0;
   assign ecchmatrix[7][77] = 0;
   assign ecchmatrix[8][77] = 1;
   assign ecchmatrix[9][77] = 0;
   assign ecchmatrix[0][78] = 0;
   assign ecchmatrix[1][78] = 0;
   assign ecchmatrix[2][78] = 1;
   assign ecchmatrix[3][78] = 0;
   assign ecchmatrix[4][78] = 0;
   assign ecchmatrix[5][78] = 1;
   assign ecchmatrix[6][78] = 0;
   assign ecchmatrix[7][78] = 0;
   assign ecchmatrix[8][78] = 0;
   assign ecchmatrix[9][78] = 1;
   assign ecchmatrix[0][79] = 0;
   assign ecchmatrix[1][79] = 0;
   assign ecchmatrix[2][79] = 1;
   assign ecchmatrix[3][79] = 0;
   assign ecchmatrix[4][79] = 0;
   assign ecchmatrix[5][79] = 0;
   assign ecchmatrix[6][79] = 1;
   assign ecchmatrix[7][79] = 1;
   assign ecchmatrix[8][79] = 0;
   assign ecchmatrix[9][79] = 0;
   assign ecchmatrix[0][80] = 0;
   assign ecchmatrix[1][80] = 0;
   assign ecchmatrix[2][80] = 1;
   assign ecchmatrix[3][80] = 0;
   assign ecchmatrix[4][80] = 0;
   assign ecchmatrix[5][80] = 0;
   assign ecchmatrix[6][80] = 1;
   assign ecchmatrix[7][80] = 0;
   assign ecchmatrix[8][80] = 1;
   assign ecchmatrix[9][80] = 0;
   assign ecchmatrix[0][81] = 0;
   assign ecchmatrix[1][81] = 0;
   assign ecchmatrix[2][81] = 1;
   assign ecchmatrix[3][81] = 0;
   assign ecchmatrix[4][81] = 0;
   assign ecchmatrix[5][81] = 0;
   assign ecchmatrix[6][81] = 1;
   assign ecchmatrix[7][81] = 0;
   assign ecchmatrix[8][81] = 0;
   assign ecchmatrix[9][81] = 1;
   assign ecchmatrix[0][82] = 0;
   assign ecchmatrix[1][82] = 0;
   assign ecchmatrix[2][82] = 1;
   assign ecchmatrix[3][82] = 0;
   assign ecchmatrix[4][82] = 0;
   assign ecchmatrix[5][82] = 0;
   assign ecchmatrix[6][82] = 0;
   assign ecchmatrix[7][82] = 1;
   assign ecchmatrix[8][82] = 1;
   assign ecchmatrix[9][82] = 0;
   assign ecchmatrix[0][83] = 0;
   assign ecchmatrix[1][83] = 0;
   assign ecchmatrix[2][83] = 1;
   assign ecchmatrix[3][83] = 0;
   assign ecchmatrix[4][83] = 0;
   assign ecchmatrix[5][83] = 0;
   assign ecchmatrix[6][83] = 0;
   assign ecchmatrix[7][83] = 1;
   assign ecchmatrix[8][83] = 0;
   assign ecchmatrix[9][83] = 1;
   assign ecchmatrix[0][84] = 0;
   assign ecchmatrix[1][84] = 0;
   assign ecchmatrix[2][84] = 1;
   assign ecchmatrix[3][84] = 0;
   assign ecchmatrix[4][84] = 0;
   assign ecchmatrix[5][84] = 0;
   assign ecchmatrix[6][84] = 0;
   assign ecchmatrix[7][84] = 0;
   assign ecchmatrix[8][84] = 1;
   assign ecchmatrix[9][84] = 1;
   assign ecchmatrix[0][85] = 0;
   assign ecchmatrix[1][85] = 0;
   assign ecchmatrix[2][85] = 0;
   assign ecchmatrix[3][85] = 1;
   assign ecchmatrix[4][85] = 1;
   assign ecchmatrix[5][85] = 1;
   assign ecchmatrix[6][85] = 0;
   assign ecchmatrix[7][85] = 0;
   assign ecchmatrix[8][85] = 0;
   assign ecchmatrix[9][85] = 0;
   assign ecchmatrix[0][86] = 0;
   assign ecchmatrix[1][86] = 0;
   assign ecchmatrix[2][86] = 0;
   assign ecchmatrix[3][86] = 1;
   assign ecchmatrix[4][86] = 1;
   assign ecchmatrix[5][86] = 0;
   assign ecchmatrix[6][86] = 1;
   assign ecchmatrix[7][86] = 0;
   assign ecchmatrix[8][86] = 0;
   assign ecchmatrix[9][86] = 0;
   assign ecchmatrix[0][87] = 0;
   assign ecchmatrix[1][87] = 0;
   assign ecchmatrix[2][87] = 0;
   assign ecchmatrix[3][87] = 1;
   assign ecchmatrix[4][87] = 1;
   assign ecchmatrix[5][87] = 0;
   assign ecchmatrix[6][87] = 0;
   assign ecchmatrix[7][87] = 1;
   assign ecchmatrix[8][87] = 0;
   assign ecchmatrix[9][87] = 0;
   assign ecchmatrix[0][88] = 0;
   assign ecchmatrix[1][88] = 0;
   assign ecchmatrix[2][88] = 0;
   assign ecchmatrix[3][88] = 1;
   assign ecchmatrix[4][88] = 1;
   assign ecchmatrix[5][88] = 0;
   assign ecchmatrix[6][88] = 0;
   assign ecchmatrix[7][88] = 0;
   assign ecchmatrix[8][88] = 1;
   assign ecchmatrix[9][88] = 0;
   assign ecchmatrix[0][89] = 0;
   assign ecchmatrix[1][89] = 0;
   assign ecchmatrix[2][89] = 0;
   assign ecchmatrix[3][89] = 1;
   assign ecchmatrix[4][89] = 1;
   assign ecchmatrix[5][89] = 0;
   assign ecchmatrix[6][89] = 0;
   assign ecchmatrix[7][89] = 0;
   assign ecchmatrix[8][89] = 0;
   assign ecchmatrix[9][89] = 1;
   assign ecchmatrix[0][90] = 0;
   assign ecchmatrix[1][90] = 0;
   assign ecchmatrix[2][90] = 0;
   assign ecchmatrix[3][90] = 1;
   assign ecchmatrix[4][90] = 0;
   assign ecchmatrix[5][90] = 1;
   assign ecchmatrix[6][90] = 1;
   assign ecchmatrix[7][90] = 0;
   assign ecchmatrix[8][90] = 0;
   assign ecchmatrix[9][90] = 0;
   assign ecchmatrix[0][91] = 0;
   assign ecchmatrix[1][91] = 0;
   assign ecchmatrix[2][91] = 0;
   assign ecchmatrix[3][91] = 1;
   assign ecchmatrix[4][91] = 0;
   assign ecchmatrix[5][91] = 1;
   assign ecchmatrix[6][91] = 0;
   assign ecchmatrix[7][91] = 1;
   assign ecchmatrix[8][91] = 0;
   assign ecchmatrix[9][91] = 0;
   assign ecchmatrix[0][92] = 0;
   assign ecchmatrix[1][92] = 0;
   assign ecchmatrix[2][92] = 0;
   assign ecchmatrix[3][92] = 1;
   assign ecchmatrix[4][92] = 0;
   assign ecchmatrix[5][92] = 1;
   assign ecchmatrix[6][92] = 0;
   assign ecchmatrix[7][92] = 0;
   assign ecchmatrix[8][92] = 1;
   assign ecchmatrix[9][92] = 0;
   assign ecchmatrix[0][93] = 0;
   assign ecchmatrix[1][93] = 0;
   assign ecchmatrix[2][93] = 0;
   assign ecchmatrix[3][93] = 1;
   assign ecchmatrix[4][93] = 0;
   assign ecchmatrix[5][93] = 1;
   assign ecchmatrix[6][93] = 0;
   assign ecchmatrix[7][93] = 0;
   assign ecchmatrix[8][93] = 0;
   assign ecchmatrix[9][93] = 1;
   assign ecchmatrix[0][94] = 0;
   assign ecchmatrix[1][94] = 0;
   assign ecchmatrix[2][94] = 0;
   assign ecchmatrix[3][94] = 1;
   assign ecchmatrix[4][94] = 0;
   assign ecchmatrix[5][94] = 0;
   assign ecchmatrix[6][94] = 1;
   assign ecchmatrix[7][94] = 1;
   assign ecchmatrix[8][94] = 0;
   assign ecchmatrix[9][94] = 0;
   assign ecchmatrix[0][95] = 0;
   assign ecchmatrix[1][95] = 0;
   assign ecchmatrix[2][95] = 0;
   assign ecchmatrix[3][95] = 1;
   assign ecchmatrix[4][95] = 0;
   assign ecchmatrix[5][95] = 0;
   assign ecchmatrix[6][95] = 1;
   assign ecchmatrix[7][95] = 0;
   assign ecchmatrix[8][95] = 1;
   assign ecchmatrix[9][95] = 0;
   assign ecchmatrix[0][96] = 0;
   assign ecchmatrix[1][96] = 0;
   assign ecchmatrix[2][96] = 0;
   assign ecchmatrix[3][96] = 1;
   assign ecchmatrix[4][96] = 0;
   assign ecchmatrix[5][96] = 0;
   assign ecchmatrix[6][96] = 1;
   assign ecchmatrix[7][96] = 0;
   assign ecchmatrix[8][96] = 0;
   assign ecchmatrix[9][96] = 1;
   assign ecchmatrix[0][97] = 0;
   assign ecchmatrix[1][97] = 0;
   assign ecchmatrix[2][97] = 0;
   assign ecchmatrix[3][97] = 1;
   assign ecchmatrix[4][97] = 0;
   assign ecchmatrix[5][97] = 0;
   assign ecchmatrix[6][97] = 0;
   assign ecchmatrix[7][97] = 1;
   assign ecchmatrix[8][97] = 1;
   assign ecchmatrix[9][97] = 0;
   assign ecchmatrix[0][98] = 0;
   assign ecchmatrix[1][98] = 0;
   assign ecchmatrix[2][98] = 0;
   assign ecchmatrix[3][98] = 1;
   assign ecchmatrix[4][98] = 0;
   assign ecchmatrix[5][98] = 0;
   assign ecchmatrix[6][98] = 0;
   assign ecchmatrix[7][98] = 1;
   assign ecchmatrix[8][98] = 0;
   assign ecchmatrix[9][98] = 1;
   assign ecchmatrix[0][99] = 0;
   assign ecchmatrix[1][99] = 0;
   assign ecchmatrix[2][99] = 0;
   assign ecchmatrix[3][99] = 1;
   assign ecchmatrix[4][99] = 0;
   assign ecchmatrix[5][99] = 0;
   assign ecchmatrix[6][99] = 0;
   assign ecchmatrix[7][99] = 0;
   assign ecchmatrix[8][99] = 1;
   assign ecchmatrix[9][99] = 1;
   assign ecchmatrix[0][100] = 0;
   assign ecchmatrix[1][100] = 0;
   assign ecchmatrix[2][100] = 0;
   assign ecchmatrix[3][100] = 0;
   assign ecchmatrix[4][100] = 1;
   assign ecchmatrix[5][100] = 1;
   assign ecchmatrix[6][100] = 1;
   assign ecchmatrix[7][100] = 0;
   assign ecchmatrix[8][100] = 0;
   assign ecchmatrix[9][100] = 0;
   assign ecchmatrix[0][101] = 0;
   assign ecchmatrix[1][101] = 0;
   assign ecchmatrix[2][101] = 0;
   assign ecchmatrix[3][101] = 0;
   assign ecchmatrix[4][101] = 1;
   assign ecchmatrix[5][101] = 1;
   assign ecchmatrix[6][101] = 0;
   assign ecchmatrix[7][101] = 1;
   assign ecchmatrix[8][101] = 0;
   assign ecchmatrix[9][101] = 0;
   assign ecchmatrix[0][102] = 0;
   assign ecchmatrix[1][102] = 0;
   assign ecchmatrix[2][102] = 0;
   assign ecchmatrix[3][102] = 0;
   assign ecchmatrix[4][102] = 1;
   assign ecchmatrix[5][102] = 1;
   assign ecchmatrix[6][102] = 0;
   assign ecchmatrix[7][102] = 0;
   assign ecchmatrix[8][102] = 1;
   assign ecchmatrix[9][102] = 0;
   assign ecchmatrix[0][103] = 0;
   assign ecchmatrix[1][103] = 0;
   assign ecchmatrix[2][103] = 0;
   assign ecchmatrix[3][103] = 0;
   assign ecchmatrix[4][103] = 1;
   assign ecchmatrix[5][103] = 1;
   assign ecchmatrix[6][103] = 0;
   assign ecchmatrix[7][103] = 0;
   assign ecchmatrix[8][103] = 0;
   assign ecchmatrix[9][103] = 1;
   assign ecchmatrix[0][104] = 0;
   assign ecchmatrix[1][104] = 0;
   assign ecchmatrix[2][104] = 0;
   assign ecchmatrix[3][104] = 0;
   assign ecchmatrix[4][104] = 1;
   assign ecchmatrix[5][104] = 0;
   assign ecchmatrix[6][104] = 1;
   assign ecchmatrix[7][104] = 1;
   assign ecchmatrix[8][104] = 0;
   assign ecchmatrix[9][104] = 0;
   assign ecchmatrix[0][105] = 0;
   assign ecchmatrix[1][105] = 0;
   assign ecchmatrix[2][105] = 0;
   assign ecchmatrix[3][105] = 0;
   assign ecchmatrix[4][105] = 1;
   assign ecchmatrix[5][105] = 0;
   assign ecchmatrix[6][105] = 1;
   assign ecchmatrix[7][105] = 0;
   assign ecchmatrix[8][105] = 1;
   assign ecchmatrix[9][105] = 0;
   assign ecchmatrix[0][106] = 0;
   assign ecchmatrix[1][106] = 0;
   assign ecchmatrix[2][106] = 0;
   assign ecchmatrix[3][106] = 0;
   assign ecchmatrix[4][106] = 1;
   assign ecchmatrix[5][106] = 0;
   assign ecchmatrix[6][106] = 1;
   assign ecchmatrix[7][106] = 0;
   assign ecchmatrix[8][106] = 0;
   assign ecchmatrix[9][106] = 1;
   assign ecchmatrix[0][107] = 0;
   assign ecchmatrix[1][107] = 0;
   assign ecchmatrix[2][107] = 0;
   assign ecchmatrix[3][107] = 0;
   assign ecchmatrix[4][107] = 1;
   assign ecchmatrix[5][107] = 0;
   assign ecchmatrix[6][107] = 0;
   assign ecchmatrix[7][107] = 1;
   assign ecchmatrix[8][107] = 1;
   assign ecchmatrix[9][107] = 0;
   assign ecchmatrix[0][108] = 0;
   assign ecchmatrix[1][108] = 0;
   assign ecchmatrix[2][108] = 0;
   assign ecchmatrix[3][108] = 0;
   assign ecchmatrix[4][108] = 1;
   assign ecchmatrix[5][108] = 0;
   assign ecchmatrix[6][108] = 0;
   assign ecchmatrix[7][108] = 1;
   assign ecchmatrix[8][108] = 0;
   assign ecchmatrix[9][108] = 1;
   assign ecchmatrix[0][109] = 0;
   assign ecchmatrix[1][109] = 0;
   assign ecchmatrix[2][109] = 0;
   assign ecchmatrix[3][109] = 0;
   assign ecchmatrix[4][109] = 1;
   assign ecchmatrix[5][109] = 0;
   assign ecchmatrix[6][109] = 0;
   assign ecchmatrix[7][109] = 0;
   assign ecchmatrix[8][109] = 1;
   assign ecchmatrix[9][109] = 1;
   assign ecchmatrix[0][110] = 0;
   assign ecchmatrix[1][110] = 0;
   assign ecchmatrix[2][110] = 0;
   assign ecchmatrix[3][110] = 0;
   assign ecchmatrix[4][110] = 0;
   assign ecchmatrix[5][110] = 1;
   assign ecchmatrix[6][110] = 1;
   assign ecchmatrix[7][110] = 1;
   assign ecchmatrix[8][110] = 0;
   assign ecchmatrix[9][110] = 0;
   assign ecchmatrix[0][111] = 0;
   assign ecchmatrix[1][111] = 0;
   assign ecchmatrix[2][111] = 0;
   assign ecchmatrix[3][111] = 0;
   assign ecchmatrix[4][111] = 0;
   assign ecchmatrix[5][111] = 1;
   assign ecchmatrix[6][111] = 1;
   assign ecchmatrix[7][111] = 0;
   assign ecchmatrix[8][111] = 1;
   assign ecchmatrix[9][111] = 0;
   assign ecchmatrix[0][112] = 0;
   assign ecchmatrix[1][112] = 0;
   assign ecchmatrix[2][112] = 0;
   assign ecchmatrix[3][112] = 0;
   assign ecchmatrix[4][112] = 0;
   assign ecchmatrix[5][112] = 1;
   assign ecchmatrix[6][112] = 1;
   assign ecchmatrix[7][112] = 0;
   assign ecchmatrix[8][112] = 0;
   assign ecchmatrix[9][112] = 1;
   assign ecchmatrix[0][113] = 0;
   assign ecchmatrix[1][113] = 0;
   assign ecchmatrix[2][113] = 0;
   assign ecchmatrix[3][113] = 0;
   assign ecchmatrix[4][113] = 0;
   assign ecchmatrix[5][113] = 1;
   assign ecchmatrix[6][113] = 0;
   assign ecchmatrix[7][113] = 1;
   assign ecchmatrix[8][113] = 1;
   assign ecchmatrix[9][113] = 0;
   assign ecchmatrix[0][114] = 0;
   assign ecchmatrix[1][114] = 0;
   assign ecchmatrix[2][114] = 0;
   assign ecchmatrix[3][114] = 0;
   assign ecchmatrix[4][114] = 0;
   assign ecchmatrix[5][114] = 1;
   assign ecchmatrix[6][114] = 0;
   assign ecchmatrix[7][114] = 1;
   assign ecchmatrix[8][114] = 0;
   assign ecchmatrix[9][114] = 1;
   assign ecchmatrix[0][115] = 0;
   assign ecchmatrix[1][115] = 0;
   assign ecchmatrix[2][115] = 0;
   assign ecchmatrix[3][115] = 0;
   assign ecchmatrix[4][115] = 0;
   assign ecchmatrix[5][115] = 1;
   assign ecchmatrix[6][115] = 0;
   assign ecchmatrix[7][115] = 0;
   assign ecchmatrix[8][115] = 1;
   assign ecchmatrix[9][115] = 1;
   assign ecchmatrix[0][116] = 0;
   assign ecchmatrix[1][116] = 0;
   assign ecchmatrix[2][116] = 0;
   assign ecchmatrix[3][116] = 0;
   assign ecchmatrix[4][116] = 0;
   assign ecchmatrix[5][116] = 0;
   assign ecchmatrix[6][116] = 1;
   assign ecchmatrix[7][116] = 1;
   assign ecchmatrix[8][116] = 1;
   assign ecchmatrix[9][116] = 0;
   assign ecchmatrix[0][117] = 0;
   assign ecchmatrix[1][117] = 0;
   assign ecchmatrix[2][117] = 0;
   assign ecchmatrix[3][117] = 0;
   assign ecchmatrix[4][117] = 0;
   assign ecchmatrix[5][117] = 0;
   assign ecchmatrix[6][117] = 1;
   assign ecchmatrix[7][117] = 1;
   assign ecchmatrix[8][117] = 0;
   assign ecchmatrix[9][117] = 1;
   assign ecchmatrix[0][118] = 0;
   assign ecchmatrix[1][118] = 0;
   assign ecchmatrix[2][118] = 0;
   assign ecchmatrix[3][118] = 0;
   assign ecchmatrix[4][118] = 0;
   assign ecchmatrix[5][118] = 0;
   assign ecchmatrix[6][118] = 1;
   assign ecchmatrix[7][118] = 0;
   assign ecchmatrix[8][118] = 1;
   assign ecchmatrix[9][118] = 1;
   assign ecchmatrix[0][119] = 0;
   assign ecchmatrix[1][119] = 0;
   assign ecchmatrix[2][119] = 0;
   assign ecchmatrix[3][119] = 0;
   assign ecchmatrix[4][119] = 0;
   assign ecchmatrix[5][119] = 0;
   assign ecchmatrix[6][119] = 0;
   assign ecchmatrix[7][119] = 1;
   assign ecchmatrix[8][119] = 1;
   assign ecchmatrix[9][119] = 1;
   assign ecchmatrix[0][120] = 1;
   assign ecchmatrix[1][120] = 1;
   assign ecchmatrix[2][120] = 1;
   assign ecchmatrix[3][120] = 1;
   assign ecchmatrix[4][120] = 1;
   assign ecchmatrix[5][120] = 0;
   assign ecchmatrix[6][120] = 0;
   assign ecchmatrix[7][120] = 0;
   assign ecchmatrix[8][120] = 0;
   assign ecchmatrix[9][120] = 0;
   assign ecchmatrix[0][121] = 1;
   assign ecchmatrix[1][121] = 1;
   assign ecchmatrix[2][121] = 1;
   assign ecchmatrix[3][121] = 1;
   assign ecchmatrix[4][121] = 0;
   assign ecchmatrix[5][121] = 1;
   assign ecchmatrix[6][121] = 0;
   assign ecchmatrix[7][121] = 0;
   assign ecchmatrix[8][121] = 0;
   assign ecchmatrix[9][121] = 0;
   assign ecchmatrix[0][122] = 1;
   assign ecchmatrix[1][122] = 1;
   assign ecchmatrix[2][122] = 1;
   assign ecchmatrix[3][122] = 1;
   assign ecchmatrix[4][122] = 0;
   assign ecchmatrix[5][122] = 0;
   assign ecchmatrix[6][122] = 1;
   assign ecchmatrix[7][122] = 0;
   assign ecchmatrix[8][122] = 0;
   assign ecchmatrix[9][122] = 0;
   assign ecchmatrix[0][123] = 1;
   assign ecchmatrix[1][123] = 1;
   assign ecchmatrix[2][123] = 1;
   assign ecchmatrix[3][123] = 1;
   assign ecchmatrix[4][123] = 0;
   assign ecchmatrix[5][123] = 0;
   assign ecchmatrix[6][123] = 0;
   assign ecchmatrix[7][123] = 1;
   assign ecchmatrix[8][123] = 0;
   assign ecchmatrix[9][123] = 0;
   assign ecchmatrix[0][124] = 1;
   assign ecchmatrix[1][124] = 1;
   assign ecchmatrix[2][124] = 1;
   assign ecchmatrix[3][124] = 1;
   assign ecchmatrix[4][124] = 0;
   assign ecchmatrix[5][124] = 0;
   assign ecchmatrix[6][124] = 0;
   assign ecchmatrix[7][124] = 0;
   assign ecchmatrix[8][124] = 1;
   assign ecchmatrix[9][124] = 0;
   assign ecchmatrix[0][125] = 1;
   assign ecchmatrix[1][125] = 1;
   assign ecchmatrix[2][125] = 1;
   assign ecchmatrix[3][125] = 1;
   assign ecchmatrix[4][125] = 0;
   assign ecchmatrix[5][125] = 0;
   assign ecchmatrix[6][125] = 0;
   assign ecchmatrix[7][125] = 0;
   assign ecchmatrix[8][125] = 0;
   assign ecchmatrix[9][125] = 1;
   assign ecchmatrix[0][126] = 1;
   assign ecchmatrix[1][126] = 1;
   assign ecchmatrix[2][126] = 1;
   assign ecchmatrix[3][126] = 0;
   assign ecchmatrix[4][126] = 1;
   assign ecchmatrix[5][126] = 1;
   assign ecchmatrix[6][126] = 0;
   assign ecchmatrix[7][126] = 0;
   assign ecchmatrix[8][126] = 0;
   assign ecchmatrix[9][126] = 0;
   assign ecchmatrix[0][127] = 1;
   assign ecchmatrix[1][127] = 1;
   assign ecchmatrix[2][127] = 1;
   assign ecchmatrix[3][127] = 0;
   assign ecchmatrix[4][127] = 1;
   assign ecchmatrix[5][127] = 0;
   assign ecchmatrix[6][127] = 1;
   assign ecchmatrix[7][127] = 0;
   assign ecchmatrix[8][127] = 0;
   assign ecchmatrix[9][127] = 0;
   assign ecchmatrix[0][128] = 1;
   assign ecchmatrix[1][128] = 1;
   assign ecchmatrix[2][128] = 1;
   assign ecchmatrix[3][128] = 0;
   assign ecchmatrix[4][128] = 1;
   assign ecchmatrix[5][128] = 0;
   assign ecchmatrix[6][128] = 0;
   assign ecchmatrix[7][128] = 1;
   assign ecchmatrix[8][128] = 0;
   assign ecchmatrix[9][128] = 0;
   assign ecchmatrix[0][129] = 1;
   assign ecchmatrix[1][129] = 1;
   assign ecchmatrix[2][129] = 1;
   assign ecchmatrix[3][129] = 0;
   assign ecchmatrix[4][129] = 1;
   assign ecchmatrix[5][129] = 0;
   assign ecchmatrix[6][129] = 0;
   assign ecchmatrix[7][129] = 0;
   assign ecchmatrix[8][129] = 1;
   assign ecchmatrix[9][129] = 0;
   assign ecchmatrix[0][130] = 1;
   assign ecchmatrix[1][130] = 1;
   assign ecchmatrix[2][130] = 1;
   assign ecchmatrix[3][130] = 0;
   assign ecchmatrix[4][130] = 1;
   assign ecchmatrix[5][130] = 0;
   assign ecchmatrix[6][130] = 0;
   assign ecchmatrix[7][130] = 0;
   assign ecchmatrix[8][130] = 0;
   assign ecchmatrix[9][130] = 1;
   assign ecchmatrix[0][131] = 1;
   assign ecchmatrix[1][131] = 1;
   assign ecchmatrix[2][131] = 1;
   assign ecchmatrix[3][131] = 0;
   assign ecchmatrix[4][131] = 0;
   assign ecchmatrix[5][131] = 1;
   assign ecchmatrix[6][131] = 1;
   assign ecchmatrix[7][131] = 0;
   assign ecchmatrix[8][131] = 0;
   assign ecchmatrix[9][131] = 0;
   assign ecchmatrix[0][132] = 1;
   assign ecchmatrix[1][132] = 1;
   assign ecchmatrix[2][132] = 1;
   assign ecchmatrix[3][132] = 0;
   assign ecchmatrix[4][132] = 0;
   assign ecchmatrix[5][132] = 1;
   assign ecchmatrix[6][132] = 0;
   assign ecchmatrix[7][132] = 1;
   assign ecchmatrix[8][132] = 0;
   assign ecchmatrix[9][132] = 0;
   assign ecchmatrix[0][133] = 1;
   assign ecchmatrix[1][133] = 1;
   assign ecchmatrix[2][133] = 1;
   assign ecchmatrix[3][133] = 0;
   assign ecchmatrix[4][133] = 0;
   assign ecchmatrix[5][133] = 1;
   assign ecchmatrix[6][133] = 0;
   assign ecchmatrix[7][133] = 0;
   assign ecchmatrix[8][133] = 1;
   assign ecchmatrix[9][133] = 0;
   assign ecchmatrix[0][134] = 1;
   assign ecchmatrix[1][134] = 1;
   assign ecchmatrix[2][134] = 1;
   assign ecchmatrix[3][134] = 0;
   assign ecchmatrix[4][134] = 0;
   assign ecchmatrix[5][134] = 1;
   assign ecchmatrix[6][134] = 0;
   assign ecchmatrix[7][134] = 0;
   assign ecchmatrix[8][134] = 0;
   assign ecchmatrix[9][134] = 1;
   assign ecchmatrix[0][135] = 1;
   assign ecchmatrix[1][135] = 1;
   assign ecchmatrix[2][135] = 1;
   assign ecchmatrix[3][135] = 0;
   assign ecchmatrix[4][135] = 0;
   assign ecchmatrix[5][135] = 0;
   assign ecchmatrix[6][135] = 1;
   assign ecchmatrix[7][135] = 1;
   assign ecchmatrix[8][135] = 0;
   assign ecchmatrix[9][135] = 0;
   assign ecchmatrix[0][136] = 1;
   assign ecchmatrix[1][136] = 1;
   assign ecchmatrix[2][136] = 1;
   assign ecchmatrix[3][136] = 0;
   assign ecchmatrix[4][136] = 0;
   assign ecchmatrix[5][136] = 0;
   assign ecchmatrix[6][136] = 1;
   assign ecchmatrix[7][136] = 0;
   assign ecchmatrix[8][136] = 1;
   assign ecchmatrix[9][136] = 0;
   assign ecchmatrix[0][137] = 1;
   assign ecchmatrix[1][137] = 1;
   assign ecchmatrix[2][137] = 1;
   assign ecchmatrix[3][137] = 0;
   assign ecchmatrix[4][137] = 0;
   assign ecchmatrix[5][137] = 0;
   assign ecchmatrix[6][137] = 1;
   assign ecchmatrix[7][137] = 0;
   assign ecchmatrix[8][137] = 0;
   assign ecchmatrix[9][137] = 1;
   assign ecchmatrix[0][138] = 1;
   assign ecchmatrix[1][138] = 1;
   assign ecchmatrix[2][138] = 1;
   assign ecchmatrix[3][138] = 0;
   assign ecchmatrix[4][138] = 0;
   assign ecchmatrix[5][138] = 0;
   assign ecchmatrix[6][138] = 0;
   assign ecchmatrix[7][138] = 1;
   assign ecchmatrix[8][138] = 1;
   assign ecchmatrix[9][138] = 0;
   assign ecchmatrix[0][139] = 1;
   assign ecchmatrix[1][139] = 1;
   assign ecchmatrix[2][139] = 1;
   assign ecchmatrix[3][139] = 0;
   assign ecchmatrix[4][139] = 0;
   assign ecchmatrix[5][139] = 0;
   assign ecchmatrix[6][139] = 0;
   assign ecchmatrix[7][139] = 1;
   assign ecchmatrix[8][139] = 0;
   assign ecchmatrix[9][139] = 1;
   assign ecchmatrix[0][140] = 1;
   assign ecchmatrix[1][140] = 1;
   assign ecchmatrix[2][140] = 1;
   assign ecchmatrix[3][140] = 0;
   assign ecchmatrix[4][140] = 0;
   assign ecchmatrix[5][140] = 0;
   assign ecchmatrix[6][140] = 0;
   assign ecchmatrix[7][140] = 0;
   assign ecchmatrix[8][140] = 1;
   assign ecchmatrix[9][140] = 1;
   assign ecchmatrix[0][141] = 1;
   assign ecchmatrix[1][141] = 1;
   assign ecchmatrix[2][141] = 0;
   assign ecchmatrix[3][141] = 1;
   assign ecchmatrix[4][141] = 1;
   assign ecchmatrix[5][141] = 1;
   assign ecchmatrix[6][141] = 0;
   assign ecchmatrix[7][141] = 0;
   assign ecchmatrix[8][141] = 0;
   assign ecchmatrix[9][141] = 0;
   assign ecchmatrix[0][142] = 1;
   assign ecchmatrix[1][142] = 1;
   assign ecchmatrix[2][142] = 0;
   assign ecchmatrix[3][142] = 1;
   assign ecchmatrix[4][142] = 1;
   assign ecchmatrix[5][142] = 0;
   assign ecchmatrix[6][142] = 1;
   assign ecchmatrix[7][142] = 0;
   assign ecchmatrix[8][142] = 0;
   assign ecchmatrix[9][142] = 0;
   assign ecchmatrix[0][143] = 1;
   assign ecchmatrix[1][143] = 1;
   assign ecchmatrix[2][143] = 0;
   assign ecchmatrix[3][143] = 1;
   assign ecchmatrix[4][143] = 1;
   assign ecchmatrix[5][143] = 0;
   assign ecchmatrix[6][143] = 0;
   assign ecchmatrix[7][143] = 1;
   assign ecchmatrix[8][143] = 0;
   assign ecchmatrix[9][143] = 0;
   assign ecchmatrix[0][144] = 1;
   assign ecchmatrix[1][144] = 1;
   assign ecchmatrix[2][144] = 0;
   assign ecchmatrix[3][144] = 1;
   assign ecchmatrix[4][144] = 1;
   assign ecchmatrix[5][144] = 0;
   assign ecchmatrix[6][144] = 0;
   assign ecchmatrix[7][144] = 0;
   assign ecchmatrix[8][144] = 1;
   assign ecchmatrix[9][144] = 0;
   assign ecchmatrix[0][145] = 1;
   assign ecchmatrix[1][145] = 1;
   assign ecchmatrix[2][145] = 0;
   assign ecchmatrix[3][145] = 1;
   assign ecchmatrix[4][145] = 1;
   assign ecchmatrix[5][145] = 0;
   assign ecchmatrix[6][145] = 0;
   assign ecchmatrix[7][145] = 0;
   assign ecchmatrix[8][145] = 0;
   assign ecchmatrix[9][145] = 1;
   assign ecchmatrix[0][146] = 1;
   assign ecchmatrix[1][146] = 1;
   assign ecchmatrix[2][146] = 0;
   assign ecchmatrix[3][146] = 1;
   assign ecchmatrix[4][146] = 0;
   assign ecchmatrix[5][146] = 1;
   assign ecchmatrix[6][146] = 1;
   assign ecchmatrix[7][146] = 0;
   assign ecchmatrix[8][146] = 0;
   assign ecchmatrix[9][146] = 0;
   assign ecchmatrix[0][147] = 1;
   assign ecchmatrix[1][147] = 1;
   assign ecchmatrix[2][147] = 0;
   assign ecchmatrix[3][147] = 1;
   assign ecchmatrix[4][147] = 0;
   assign ecchmatrix[5][147] = 1;
   assign ecchmatrix[6][147] = 0;
   assign ecchmatrix[7][147] = 1;
   assign ecchmatrix[8][147] = 0;
   assign ecchmatrix[9][147] = 0;
   assign ecchmatrix[0][148] = 1;
   assign ecchmatrix[1][148] = 1;
   assign ecchmatrix[2][148] = 0;
   assign ecchmatrix[3][148] = 1;
   assign ecchmatrix[4][148] = 0;
   assign ecchmatrix[5][148] = 1;
   assign ecchmatrix[6][148] = 0;
   assign ecchmatrix[7][148] = 0;
   assign ecchmatrix[8][148] = 1;
   assign ecchmatrix[9][148] = 0;
   assign ecchmatrix[0][149] = 1;
   assign ecchmatrix[1][149] = 1;
   assign ecchmatrix[2][149] = 0;
   assign ecchmatrix[3][149] = 1;
   assign ecchmatrix[4][149] = 0;
   assign ecchmatrix[5][149] = 1;
   assign ecchmatrix[6][149] = 0;
   assign ecchmatrix[7][149] = 0;
   assign ecchmatrix[8][149] = 0;
   assign ecchmatrix[9][149] = 1;
   assign ecchmatrix[0][150] = 1;
   assign ecchmatrix[1][150] = 1;
   assign ecchmatrix[2][150] = 0;
   assign ecchmatrix[3][150] = 1;
   assign ecchmatrix[4][150] = 0;
   assign ecchmatrix[5][150] = 0;
   assign ecchmatrix[6][150] = 1;
   assign ecchmatrix[7][150] = 1;
   assign ecchmatrix[8][150] = 0;
   assign ecchmatrix[9][150] = 0;
   assign ecchmatrix[0][151] = 1;
   assign ecchmatrix[1][151] = 1;
   assign ecchmatrix[2][151] = 0;
   assign ecchmatrix[3][151] = 1;
   assign ecchmatrix[4][151] = 0;
   assign ecchmatrix[5][151] = 0;
   assign ecchmatrix[6][151] = 1;
   assign ecchmatrix[7][151] = 0;
   assign ecchmatrix[8][151] = 1;
   assign ecchmatrix[9][151] = 0;
   assign ecchmatrix[0][152] = 1;
   assign ecchmatrix[1][152] = 1;
   assign ecchmatrix[2][152] = 0;
   assign ecchmatrix[3][152] = 1;
   assign ecchmatrix[4][152] = 0;
   assign ecchmatrix[5][152] = 0;
   assign ecchmatrix[6][152] = 1;
   assign ecchmatrix[7][152] = 0;
   assign ecchmatrix[8][152] = 0;
   assign ecchmatrix[9][152] = 1;
   assign ecchmatrix[0][153] = 1;
   assign ecchmatrix[1][153] = 1;
   assign ecchmatrix[2][153] = 0;
   assign ecchmatrix[3][153] = 1;
   assign ecchmatrix[4][153] = 0;
   assign ecchmatrix[5][153] = 0;
   assign ecchmatrix[6][153] = 0;
   assign ecchmatrix[7][153] = 1;
   assign ecchmatrix[8][153] = 1;
   assign ecchmatrix[9][153] = 0;
   assign ecchmatrix[0][154] = 1;
   assign ecchmatrix[1][154] = 1;
   assign ecchmatrix[2][154] = 0;
   assign ecchmatrix[3][154] = 1;
   assign ecchmatrix[4][154] = 0;
   assign ecchmatrix[5][154] = 0;
   assign ecchmatrix[6][154] = 0;
   assign ecchmatrix[7][154] = 1;
   assign ecchmatrix[8][154] = 0;
   assign ecchmatrix[9][154] = 1;
   assign ecchmatrix[0][155] = 1;
   assign ecchmatrix[1][155] = 1;
   assign ecchmatrix[2][155] = 0;
   assign ecchmatrix[3][155] = 1;
   assign ecchmatrix[4][155] = 0;
   assign ecchmatrix[5][155] = 0;
   assign ecchmatrix[6][155] = 0;
   assign ecchmatrix[7][155] = 0;
   assign ecchmatrix[8][155] = 1;
   assign ecchmatrix[9][155] = 1;
   assign ecchmatrix[0][156] = 1;
   assign ecchmatrix[1][156] = 1;
   assign ecchmatrix[2][156] = 0;
   assign ecchmatrix[3][156] = 0;
   assign ecchmatrix[4][156] = 1;
   assign ecchmatrix[5][156] = 1;
   assign ecchmatrix[6][156] = 1;
   assign ecchmatrix[7][156] = 0;
   assign ecchmatrix[8][156] = 0;
   assign ecchmatrix[9][156] = 0;
   assign ecchmatrix[0][157] = 1;
   assign ecchmatrix[1][157] = 1;
   assign ecchmatrix[2][157] = 0;
   assign ecchmatrix[3][157] = 0;
   assign ecchmatrix[4][157] = 1;
   assign ecchmatrix[5][157] = 1;
   assign ecchmatrix[6][157] = 0;
   assign ecchmatrix[7][157] = 1;
   assign ecchmatrix[8][157] = 0;
   assign ecchmatrix[9][157] = 0;
   assign ecchmatrix[0][158] = 1;
   assign ecchmatrix[1][158] = 1;
   assign ecchmatrix[2][158] = 0;
   assign ecchmatrix[3][158] = 0;
   assign ecchmatrix[4][158] = 1;
   assign ecchmatrix[5][158] = 1;
   assign ecchmatrix[6][158] = 0;
   assign ecchmatrix[7][158] = 0;
   assign ecchmatrix[8][158] = 1;
   assign ecchmatrix[9][158] = 0;
   assign ecchmatrix[0][159] = 1;
   assign ecchmatrix[1][159] = 1;
   assign ecchmatrix[2][159] = 0;
   assign ecchmatrix[3][159] = 0;
   assign ecchmatrix[4][159] = 1;
   assign ecchmatrix[5][159] = 1;
   assign ecchmatrix[6][159] = 0;
   assign ecchmatrix[7][159] = 0;
   assign ecchmatrix[8][159] = 0;
   assign ecchmatrix[9][159] = 1;
   assign ecchmatrix[0][160] = 1;
   assign ecchmatrix[1][160] = 1;
   assign ecchmatrix[2][160] = 0;
   assign ecchmatrix[3][160] = 0;
   assign ecchmatrix[4][160] = 1;
   assign ecchmatrix[5][160] = 0;
   assign ecchmatrix[6][160] = 1;
   assign ecchmatrix[7][160] = 1;
   assign ecchmatrix[8][160] = 0;
   assign ecchmatrix[9][160] = 0;
   assign ecchmatrix[0][161] = 1;
   assign ecchmatrix[1][161] = 1;
   assign ecchmatrix[2][161] = 0;
   assign ecchmatrix[3][161] = 0;
   assign ecchmatrix[4][161] = 1;
   assign ecchmatrix[5][161] = 0;
   assign ecchmatrix[6][161] = 1;
   assign ecchmatrix[7][161] = 0;
   assign ecchmatrix[8][161] = 1;
   assign ecchmatrix[9][161] = 0;
   assign ecchmatrix[0][162] = 1;
   assign ecchmatrix[1][162] = 1;
   assign ecchmatrix[2][162] = 0;
   assign ecchmatrix[3][162] = 0;
   assign ecchmatrix[4][162] = 1;
   assign ecchmatrix[5][162] = 0;
   assign ecchmatrix[6][162] = 1;
   assign ecchmatrix[7][162] = 0;
   assign ecchmatrix[8][162] = 0;
   assign ecchmatrix[9][162] = 1;
   assign ecchmatrix[0][163] = 1;
   assign ecchmatrix[1][163] = 1;
   assign ecchmatrix[2][163] = 0;
   assign ecchmatrix[3][163] = 0;
   assign ecchmatrix[4][163] = 1;
   assign ecchmatrix[5][163] = 0;
   assign ecchmatrix[6][163] = 0;
   assign ecchmatrix[7][163] = 1;
   assign ecchmatrix[8][163] = 1;
   assign ecchmatrix[9][163] = 0;
   assign ecchmatrix[0][164] = 1;
   assign ecchmatrix[1][164] = 1;
   assign ecchmatrix[2][164] = 0;
   assign ecchmatrix[3][164] = 0;
   assign ecchmatrix[4][164] = 1;
   assign ecchmatrix[5][164] = 0;
   assign ecchmatrix[6][164] = 0;
   assign ecchmatrix[7][164] = 1;
   assign ecchmatrix[8][164] = 0;
   assign ecchmatrix[9][164] = 1;
   assign ecchmatrix[0][165] = 1;
   assign ecchmatrix[1][165] = 1;
   assign ecchmatrix[2][165] = 0;
   assign ecchmatrix[3][165] = 0;
   assign ecchmatrix[4][165] = 1;
   assign ecchmatrix[5][165] = 0;
   assign ecchmatrix[6][165] = 0;
   assign ecchmatrix[7][165] = 0;
   assign ecchmatrix[8][165] = 1;
   assign ecchmatrix[9][165] = 1;
   assign ecchmatrix[0][166] = 1;
   assign ecchmatrix[1][166] = 1;
   assign ecchmatrix[2][166] = 0;
   assign ecchmatrix[3][166] = 0;
   assign ecchmatrix[4][166] = 0;
   assign ecchmatrix[5][166] = 1;
   assign ecchmatrix[6][166] = 1;
   assign ecchmatrix[7][166] = 1;
   assign ecchmatrix[8][166] = 0;
   assign ecchmatrix[9][166] = 0;
   assign ecchmatrix[0][167] = 1;
   assign ecchmatrix[1][167] = 1;
   assign ecchmatrix[2][167] = 0;
   assign ecchmatrix[3][167] = 0;
   assign ecchmatrix[4][167] = 0;
   assign ecchmatrix[5][167] = 1;
   assign ecchmatrix[6][167] = 1;
   assign ecchmatrix[7][167] = 0;
   assign ecchmatrix[8][167] = 1;
   assign ecchmatrix[9][167] = 0;
   assign ecchmatrix[0][168] = 1;
   assign ecchmatrix[1][168] = 1;
   assign ecchmatrix[2][168] = 0;
   assign ecchmatrix[3][168] = 0;
   assign ecchmatrix[4][168] = 0;
   assign ecchmatrix[5][168] = 1;
   assign ecchmatrix[6][168] = 1;
   assign ecchmatrix[7][168] = 0;
   assign ecchmatrix[8][168] = 0;
   assign ecchmatrix[9][168] = 1;
   assign ecchmatrix[0][169] = 1;
   assign ecchmatrix[1][169] = 1;
   assign ecchmatrix[2][169] = 0;
   assign ecchmatrix[3][169] = 0;
   assign ecchmatrix[4][169] = 0;
   assign ecchmatrix[5][169] = 1;
   assign ecchmatrix[6][169] = 0;
   assign ecchmatrix[7][169] = 1;
   assign ecchmatrix[8][169] = 1;
   assign ecchmatrix[9][169] = 0;
   assign ecchmatrix[0][170] = 1;
   assign ecchmatrix[1][170] = 1;
   assign ecchmatrix[2][170] = 0;
   assign ecchmatrix[3][170] = 0;
   assign ecchmatrix[4][170] = 0;
   assign ecchmatrix[5][170] = 1;
   assign ecchmatrix[6][170] = 0;
   assign ecchmatrix[7][170] = 1;
   assign ecchmatrix[8][170] = 0;
   assign ecchmatrix[9][170] = 1;
   assign ecchmatrix[0][171] = 1;
   assign ecchmatrix[1][171] = 1;
   assign ecchmatrix[2][171] = 0;
   assign ecchmatrix[3][171] = 0;
   assign ecchmatrix[4][171] = 0;
   assign ecchmatrix[5][171] = 1;
   assign ecchmatrix[6][171] = 0;
   assign ecchmatrix[7][171] = 0;
   assign ecchmatrix[8][171] = 1;
   assign ecchmatrix[9][171] = 1;
   assign ecchmatrix[0][172] = 1;
   assign ecchmatrix[1][172] = 1;
   assign ecchmatrix[2][172] = 0;
   assign ecchmatrix[3][172] = 0;
   assign ecchmatrix[4][172] = 0;
   assign ecchmatrix[5][172] = 0;
   assign ecchmatrix[6][172] = 1;
   assign ecchmatrix[7][172] = 1;
   assign ecchmatrix[8][172] = 1;
   assign ecchmatrix[9][172] = 0;
   assign ecchmatrix[0][173] = 1;
   assign ecchmatrix[1][173] = 1;
   assign ecchmatrix[2][173] = 0;
   assign ecchmatrix[3][173] = 0;
   assign ecchmatrix[4][173] = 0;
   assign ecchmatrix[5][173] = 0;
   assign ecchmatrix[6][173] = 1;
   assign ecchmatrix[7][173] = 1;
   assign ecchmatrix[8][173] = 0;
   assign ecchmatrix[9][173] = 1;
   assign ecchmatrix[0][174] = 1;
   assign ecchmatrix[1][174] = 1;
   assign ecchmatrix[2][174] = 0;
   assign ecchmatrix[3][174] = 0;
   assign ecchmatrix[4][174] = 0;
   assign ecchmatrix[5][174] = 0;
   assign ecchmatrix[6][174] = 1;
   assign ecchmatrix[7][174] = 0;
   assign ecchmatrix[8][174] = 1;
   assign ecchmatrix[9][174] = 1;
   assign ecchmatrix[0][175] = 1;
   assign ecchmatrix[1][175] = 1;
   assign ecchmatrix[2][175] = 0;
   assign ecchmatrix[3][175] = 0;
   assign ecchmatrix[4][175] = 0;
   assign ecchmatrix[5][175] = 0;
   assign ecchmatrix[6][175] = 0;
   assign ecchmatrix[7][175] = 1;
   assign ecchmatrix[8][175] = 1;
   assign ecchmatrix[9][175] = 1;
   assign ecchmatrix[0][176] = 1;
   assign ecchmatrix[1][176] = 0;
   assign ecchmatrix[2][176] = 1;
   assign ecchmatrix[3][176] = 1;
   assign ecchmatrix[4][176] = 1;
   assign ecchmatrix[5][176] = 1;
   assign ecchmatrix[6][176] = 0;
   assign ecchmatrix[7][176] = 0;
   assign ecchmatrix[8][176] = 0;
   assign ecchmatrix[9][176] = 0;
   assign ecchmatrix[0][177] = 1;
   assign ecchmatrix[1][177] = 0;
   assign ecchmatrix[2][177] = 1;
   assign ecchmatrix[3][177] = 1;
   assign ecchmatrix[4][177] = 1;
   assign ecchmatrix[5][177] = 0;
   assign ecchmatrix[6][177] = 1;
   assign ecchmatrix[7][177] = 0;
   assign ecchmatrix[8][177] = 0;
   assign ecchmatrix[9][177] = 0;
   assign ecchmatrix[0][178] = 1;
   assign ecchmatrix[1][178] = 0;
   assign ecchmatrix[2][178] = 1;
   assign ecchmatrix[3][178] = 1;
   assign ecchmatrix[4][178] = 1;
   assign ecchmatrix[5][178] = 0;
   assign ecchmatrix[6][178] = 0;
   assign ecchmatrix[7][178] = 1;
   assign ecchmatrix[8][178] = 0;
   assign ecchmatrix[9][178] = 0;
   assign ecchmatrix[0][179] = 1;
   assign ecchmatrix[1][179] = 0;
   assign ecchmatrix[2][179] = 1;
   assign ecchmatrix[3][179] = 1;
   assign ecchmatrix[4][179] = 1;
   assign ecchmatrix[5][179] = 0;
   assign ecchmatrix[6][179] = 0;
   assign ecchmatrix[7][179] = 0;
   assign ecchmatrix[8][179] = 1;
   assign ecchmatrix[9][179] = 0;
   assign ecchmatrix[0][180] = 1;
   assign ecchmatrix[1][180] = 0;
   assign ecchmatrix[2][180] = 1;
   assign ecchmatrix[3][180] = 1;
   assign ecchmatrix[4][180] = 1;
   assign ecchmatrix[5][180] = 0;
   assign ecchmatrix[6][180] = 0;
   assign ecchmatrix[7][180] = 0;
   assign ecchmatrix[8][180] = 0;
   assign ecchmatrix[9][180] = 1;
   assign ecchmatrix[0][181] = 1;
   assign ecchmatrix[1][181] = 0;
   assign ecchmatrix[2][181] = 1;
   assign ecchmatrix[3][181] = 1;
   assign ecchmatrix[4][181] = 0;
   assign ecchmatrix[5][181] = 1;
   assign ecchmatrix[6][181] = 1;
   assign ecchmatrix[7][181] = 0;
   assign ecchmatrix[8][181] = 0;
   assign ecchmatrix[9][181] = 0;
   assign ecchmatrix[0][182] = 1;
   assign ecchmatrix[1][182] = 0;
   assign ecchmatrix[2][182] = 1;
   assign ecchmatrix[3][182] = 1;
   assign ecchmatrix[4][182] = 0;
   assign ecchmatrix[5][182] = 1;
   assign ecchmatrix[6][182] = 0;
   assign ecchmatrix[7][182] = 1;
   assign ecchmatrix[8][182] = 0;
   assign ecchmatrix[9][182] = 0;
   assign ecchmatrix[0][183] = 1;
   assign ecchmatrix[1][183] = 0;
   assign ecchmatrix[2][183] = 1;
   assign ecchmatrix[3][183] = 1;
   assign ecchmatrix[4][183] = 0;
   assign ecchmatrix[5][183] = 1;
   assign ecchmatrix[6][183] = 0;
   assign ecchmatrix[7][183] = 0;
   assign ecchmatrix[8][183] = 1;
   assign ecchmatrix[9][183] = 0;
   assign ecchmatrix[0][184] = 1;
   assign ecchmatrix[1][184] = 0;
   assign ecchmatrix[2][184] = 1;
   assign ecchmatrix[3][184] = 1;
   assign ecchmatrix[4][184] = 0;
   assign ecchmatrix[5][184] = 1;
   assign ecchmatrix[6][184] = 0;
   assign ecchmatrix[7][184] = 0;
   assign ecchmatrix[8][184] = 0;
   assign ecchmatrix[9][184] = 1;
   assign ecchmatrix[0][185] = 1;
   assign ecchmatrix[1][185] = 0;
   assign ecchmatrix[2][185] = 1;
   assign ecchmatrix[3][185] = 1;
   assign ecchmatrix[4][185] = 0;
   assign ecchmatrix[5][185] = 0;
   assign ecchmatrix[6][185] = 1;
   assign ecchmatrix[7][185] = 1;
   assign ecchmatrix[8][185] = 0;
   assign ecchmatrix[9][185] = 0;
   assign ecchmatrix[0][186] = 1;
   assign ecchmatrix[1][186] = 0;
   assign ecchmatrix[2][186] = 1;
   assign ecchmatrix[3][186] = 1;
   assign ecchmatrix[4][186] = 0;
   assign ecchmatrix[5][186] = 0;
   assign ecchmatrix[6][186] = 1;
   assign ecchmatrix[7][186] = 0;
   assign ecchmatrix[8][186] = 1;
   assign ecchmatrix[9][186] = 0;
   assign ecchmatrix[0][187] = 1;
   assign ecchmatrix[1][187] = 0;
   assign ecchmatrix[2][187] = 1;
   assign ecchmatrix[3][187] = 1;
   assign ecchmatrix[4][187] = 0;
   assign ecchmatrix[5][187] = 0;
   assign ecchmatrix[6][187] = 1;
   assign ecchmatrix[7][187] = 0;
   assign ecchmatrix[8][187] = 0;
   assign ecchmatrix[9][187] = 1;
   assign ecchmatrix[0][188] = 1;
   assign ecchmatrix[1][188] = 0;
   assign ecchmatrix[2][188] = 1;
   assign ecchmatrix[3][188] = 1;
   assign ecchmatrix[4][188] = 0;
   assign ecchmatrix[5][188] = 0;
   assign ecchmatrix[6][188] = 0;
   assign ecchmatrix[7][188] = 1;
   assign ecchmatrix[8][188] = 1;
   assign ecchmatrix[9][188] = 0;
   assign ecchmatrix[0][189] = 1;
   assign ecchmatrix[1][189] = 0;
   assign ecchmatrix[2][189] = 1;
   assign ecchmatrix[3][189] = 1;
   assign ecchmatrix[4][189] = 0;
   assign ecchmatrix[5][189] = 0;
   assign ecchmatrix[6][189] = 0;
   assign ecchmatrix[7][189] = 1;
   assign ecchmatrix[8][189] = 0;
   assign ecchmatrix[9][189] = 1;
   assign ecchmatrix[0][190] = 1;
   assign ecchmatrix[1][190] = 0;
   assign ecchmatrix[2][190] = 1;
   assign ecchmatrix[3][190] = 1;
   assign ecchmatrix[4][190] = 0;
   assign ecchmatrix[5][190] = 0;
   assign ecchmatrix[6][190] = 0;
   assign ecchmatrix[7][190] = 0;
   assign ecchmatrix[8][190] = 1;
   assign ecchmatrix[9][190] = 1;
   assign ecchmatrix[0][191] = 1;
   assign ecchmatrix[1][191] = 0;
   assign ecchmatrix[2][191] = 1;
   assign ecchmatrix[3][191] = 0;
   assign ecchmatrix[4][191] = 1;
   assign ecchmatrix[5][191] = 1;
   assign ecchmatrix[6][191] = 1;
   assign ecchmatrix[7][191] = 0;
   assign ecchmatrix[8][191] = 0;
   assign ecchmatrix[9][191] = 0;
   assign ecchmatrix[0][192] = 1;
   assign ecchmatrix[1][192] = 0;
   assign ecchmatrix[2][192] = 1;
   assign ecchmatrix[3][192] = 0;
   assign ecchmatrix[4][192] = 1;
   assign ecchmatrix[5][192] = 1;
   assign ecchmatrix[6][192] = 0;
   assign ecchmatrix[7][192] = 1;
   assign ecchmatrix[8][192] = 0;
   assign ecchmatrix[9][192] = 0;
   assign ecchmatrix[0][193] = 1;
   assign ecchmatrix[1][193] = 0;
   assign ecchmatrix[2][193] = 1;
   assign ecchmatrix[3][193] = 0;
   assign ecchmatrix[4][193] = 1;
   assign ecchmatrix[5][193] = 1;
   assign ecchmatrix[6][193] = 0;
   assign ecchmatrix[7][193] = 0;
   assign ecchmatrix[8][193] = 1;
   assign ecchmatrix[9][193] = 0;
   assign ecchmatrix[0][194] = 1;
   assign ecchmatrix[1][194] = 0;
   assign ecchmatrix[2][194] = 1;
   assign ecchmatrix[3][194] = 0;
   assign ecchmatrix[4][194] = 1;
   assign ecchmatrix[5][194] = 1;
   assign ecchmatrix[6][194] = 0;
   assign ecchmatrix[7][194] = 0;
   assign ecchmatrix[8][194] = 0;
   assign ecchmatrix[9][194] = 1;
   assign ecchmatrix[0][195] = 1;
   assign ecchmatrix[1][195] = 0;
   assign ecchmatrix[2][195] = 1;
   assign ecchmatrix[3][195] = 0;
   assign ecchmatrix[4][195] = 1;
   assign ecchmatrix[5][195] = 0;
   assign ecchmatrix[6][195] = 1;
   assign ecchmatrix[7][195] = 1;
   assign ecchmatrix[8][195] = 0;
   assign ecchmatrix[9][195] = 0;
   assign ecchmatrix[0][196] = 1;
   assign ecchmatrix[1][196] = 0;
   assign ecchmatrix[2][196] = 1;
   assign ecchmatrix[3][196] = 0;
   assign ecchmatrix[4][196] = 1;
   assign ecchmatrix[5][196] = 0;
   assign ecchmatrix[6][196] = 1;
   assign ecchmatrix[7][196] = 0;
   assign ecchmatrix[8][196] = 1;
   assign ecchmatrix[9][196] = 0;
   assign ecchmatrix[0][197] = 1;
   assign ecchmatrix[1][197] = 0;
   assign ecchmatrix[2][197] = 1;
   assign ecchmatrix[3][197] = 0;
   assign ecchmatrix[4][197] = 1;
   assign ecchmatrix[5][197] = 0;
   assign ecchmatrix[6][197] = 1;
   assign ecchmatrix[7][197] = 0;
   assign ecchmatrix[8][197] = 0;
   assign ecchmatrix[9][197] = 1;
   assign ecchmatrix[0][198] = 1;
   assign ecchmatrix[1][198] = 0;
   assign ecchmatrix[2][198] = 1;
   assign ecchmatrix[3][198] = 0;
   assign ecchmatrix[4][198] = 1;
   assign ecchmatrix[5][198] = 0;
   assign ecchmatrix[6][198] = 0;
   assign ecchmatrix[7][198] = 1;
   assign ecchmatrix[8][198] = 1;
   assign ecchmatrix[9][198] = 0;
   assign ecchmatrix[0][199] = 1;
   assign ecchmatrix[1][199] = 0;
   assign ecchmatrix[2][199] = 1;
   assign ecchmatrix[3][199] = 0;
   assign ecchmatrix[4][199] = 1;
   assign ecchmatrix[5][199] = 0;
   assign ecchmatrix[6][199] = 0;
   assign ecchmatrix[7][199] = 1;
   assign ecchmatrix[8][199] = 0;
   assign ecchmatrix[9][199] = 1;
   assign ecchmatrix[0][200] = 1;
   assign ecchmatrix[1][200] = 0;
   assign ecchmatrix[2][200] = 1;
   assign ecchmatrix[3][200] = 0;
   assign ecchmatrix[4][200] = 1;
   assign ecchmatrix[5][200] = 0;
   assign ecchmatrix[6][200] = 0;
   assign ecchmatrix[7][200] = 0;
   assign ecchmatrix[8][200] = 1;
   assign ecchmatrix[9][200] = 1;
   assign ecchmatrix[0][201] = 1;
   assign ecchmatrix[1][201] = 0;
   assign ecchmatrix[2][201] = 1;
   assign ecchmatrix[3][201] = 0;
   assign ecchmatrix[4][201] = 0;
   assign ecchmatrix[5][201] = 1;
   assign ecchmatrix[6][201] = 1;
   assign ecchmatrix[7][201] = 1;
   assign ecchmatrix[8][201] = 0;
   assign ecchmatrix[9][201] = 0;
   assign ecchmatrix[0][202] = 1;
   assign ecchmatrix[1][202] = 0;
   assign ecchmatrix[2][202] = 1;
   assign ecchmatrix[3][202] = 0;
   assign ecchmatrix[4][202] = 0;
   assign ecchmatrix[5][202] = 1;
   assign ecchmatrix[6][202] = 1;
   assign ecchmatrix[7][202] = 0;
   assign ecchmatrix[8][202] = 1;
   assign ecchmatrix[9][202] = 0;
   assign ecchmatrix[0][203] = 1;
   assign ecchmatrix[1][203] = 0;
   assign ecchmatrix[2][203] = 1;
   assign ecchmatrix[3][203] = 0;
   assign ecchmatrix[4][203] = 0;
   assign ecchmatrix[5][203] = 1;
   assign ecchmatrix[6][203] = 1;
   assign ecchmatrix[7][203] = 0;
   assign ecchmatrix[8][203] = 0;
   assign ecchmatrix[9][203] = 1;
   assign ecchmatrix[0][204] = 1;
   assign ecchmatrix[1][204] = 0;
   assign ecchmatrix[2][204] = 1;
   assign ecchmatrix[3][204] = 0;
   assign ecchmatrix[4][204] = 0;
   assign ecchmatrix[5][204] = 1;
   assign ecchmatrix[6][204] = 0;
   assign ecchmatrix[7][204] = 1;
   assign ecchmatrix[8][204] = 1;
   assign ecchmatrix[9][204] = 0;
   assign ecchmatrix[0][205] = 1;
   assign ecchmatrix[1][205] = 0;
   assign ecchmatrix[2][205] = 1;
   assign ecchmatrix[3][205] = 0;
   assign ecchmatrix[4][205] = 0;
   assign ecchmatrix[5][205] = 1;
   assign ecchmatrix[6][205] = 0;
   assign ecchmatrix[7][205] = 1;
   assign ecchmatrix[8][205] = 0;
   assign ecchmatrix[9][205] = 1;
   assign ecchmatrix[0][206] = 1;
   assign ecchmatrix[1][206] = 0;
   assign ecchmatrix[2][206] = 1;
   assign ecchmatrix[3][206] = 0;
   assign ecchmatrix[4][206] = 0;
   assign ecchmatrix[5][206] = 1;
   assign ecchmatrix[6][206] = 0;
   assign ecchmatrix[7][206] = 0;
   assign ecchmatrix[8][206] = 1;
   assign ecchmatrix[9][206] = 1;
   assign ecchmatrix[0][207] = 1;
   assign ecchmatrix[1][207] = 0;
   assign ecchmatrix[2][207] = 1;
   assign ecchmatrix[3][207] = 0;
   assign ecchmatrix[4][207] = 0;
   assign ecchmatrix[5][207] = 0;
   assign ecchmatrix[6][207] = 1;
   assign ecchmatrix[7][207] = 1;
   assign ecchmatrix[8][207] = 1;
   assign ecchmatrix[9][207] = 0;
   assign ecchmatrix[0][208] = 1;
   assign ecchmatrix[1][208] = 0;
   assign ecchmatrix[2][208] = 1;
   assign ecchmatrix[3][208] = 0;
   assign ecchmatrix[4][208] = 0;
   assign ecchmatrix[5][208] = 0;
   assign ecchmatrix[6][208] = 1;
   assign ecchmatrix[7][208] = 1;
   assign ecchmatrix[8][208] = 0;
   assign ecchmatrix[9][208] = 1;
   assign ecchmatrix[0][209] = 1;
   assign ecchmatrix[1][209] = 0;
   assign ecchmatrix[2][209] = 1;
   assign ecchmatrix[3][209] = 0;
   assign ecchmatrix[4][209] = 0;
   assign ecchmatrix[5][209] = 0;
   assign ecchmatrix[6][209] = 1;
   assign ecchmatrix[7][209] = 0;
   assign ecchmatrix[8][209] = 1;
   assign ecchmatrix[9][209] = 1;
   assign ecchmatrix[0][210] = 1;
   assign ecchmatrix[1][210] = 0;
   assign ecchmatrix[2][210] = 1;
   assign ecchmatrix[3][210] = 0;
   assign ecchmatrix[4][210] = 0;
   assign ecchmatrix[5][210] = 0;
   assign ecchmatrix[6][210] = 0;
   assign ecchmatrix[7][210] = 1;
   assign ecchmatrix[8][210] = 1;
   assign ecchmatrix[9][210] = 1;
   assign ecchmatrix[0][211] = 1;
   assign ecchmatrix[1][211] = 0;
   assign ecchmatrix[2][211] = 0;
   assign ecchmatrix[3][211] = 1;
   assign ecchmatrix[4][211] = 1;
   assign ecchmatrix[5][211] = 1;
   assign ecchmatrix[6][211] = 1;
   assign ecchmatrix[7][211] = 0;
   assign ecchmatrix[8][211] = 0;
   assign ecchmatrix[9][211] = 0;
   assign ecchmatrix[0][212] = 1;
   assign ecchmatrix[1][212] = 0;
   assign ecchmatrix[2][212] = 0;
   assign ecchmatrix[3][212] = 1;
   assign ecchmatrix[4][212] = 1;
   assign ecchmatrix[5][212] = 1;
   assign ecchmatrix[6][212] = 0;
   assign ecchmatrix[7][212] = 1;
   assign ecchmatrix[8][212] = 0;
   assign ecchmatrix[9][212] = 0;
   assign ecchmatrix[0][213] = 1;
   assign ecchmatrix[1][213] = 0;
   assign ecchmatrix[2][213] = 0;
   assign ecchmatrix[3][213] = 1;
   assign ecchmatrix[4][213] = 1;
   assign ecchmatrix[5][213] = 1;
   assign ecchmatrix[6][213] = 0;
   assign ecchmatrix[7][213] = 0;
   assign ecchmatrix[8][213] = 1;
   assign ecchmatrix[9][213] = 0;
   assign ecchmatrix[0][214] = 1;
   assign ecchmatrix[1][214] = 0;
   assign ecchmatrix[2][214] = 0;
   assign ecchmatrix[3][214] = 1;
   assign ecchmatrix[4][214] = 1;
   assign ecchmatrix[5][214] = 1;
   assign ecchmatrix[6][214] = 0;
   assign ecchmatrix[7][214] = 0;
   assign ecchmatrix[8][214] = 0;
   assign ecchmatrix[9][214] = 1;
   assign ecchmatrix[0][215] = 1;
   assign ecchmatrix[1][215] = 0;
   assign ecchmatrix[2][215] = 0;
   assign ecchmatrix[3][215] = 1;
   assign ecchmatrix[4][215] = 1;
   assign ecchmatrix[5][215] = 0;
   assign ecchmatrix[6][215] = 1;
   assign ecchmatrix[7][215] = 1;
   assign ecchmatrix[8][215] = 0;
   assign ecchmatrix[9][215] = 0;
   assign ecchmatrix[0][216] = 1;
   assign ecchmatrix[1][216] = 0;
   assign ecchmatrix[2][216] = 0;
   assign ecchmatrix[3][216] = 1;
   assign ecchmatrix[4][216] = 1;
   assign ecchmatrix[5][216] = 0;
   assign ecchmatrix[6][216] = 1;
   assign ecchmatrix[7][216] = 0;
   assign ecchmatrix[8][216] = 1;
   assign ecchmatrix[9][216] = 0;
   assign ecchmatrix[0][217] = 1;
   assign ecchmatrix[1][217] = 0;
   assign ecchmatrix[2][217] = 0;
   assign ecchmatrix[3][217] = 1;
   assign ecchmatrix[4][217] = 1;
   assign ecchmatrix[5][217] = 0;
   assign ecchmatrix[6][217] = 1;
   assign ecchmatrix[7][217] = 0;
   assign ecchmatrix[8][217] = 0;
   assign ecchmatrix[9][217] = 1;
   assign ecchmatrix[0][218] = 1;
   assign ecchmatrix[1][218] = 0;
   assign ecchmatrix[2][218] = 0;
   assign ecchmatrix[3][218] = 1;
   assign ecchmatrix[4][218] = 1;
   assign ecchmatrix[5][218] = 0;
   assign ecchmatrix[6][218] = 0;
   assign ecchmatrix[7][218] = 1;
   assign ecchmatrix[8][218] = 1;
   assign ecchmatrix[9][218] = 0;
   assign ecchmatrix[0][219] = 1;
   assign ecchmatrix[1][219] = 0;
   assign ecchmatrix[2][219] = 0;
   assign ecchmatrix[3][219] = 1;
   assign ecchmatrix[4][219] = 1;
   assign ecchmatrix[5][219] = 0;
   assign ecchmatrix[6][219] = 0;
   assign ecchmatrix[7][219] = 1;
   assign ecchmatrix[8][219] = 0;
   assign ecchmatrix[9][219] = 1;
   assign ecchmatrix[0][220] = 1;
   assign ecchmatrix[1][220] = 0;
   assign ecchmatrix[2][220] = 0;
   assign ecchmatrix[3][220] = 1;
   assign ecchmatrix[4][220] = 1;
   assign ecchmatrix[5][220] = 0;
   assign ecchmatrix[6][220] = 0;
   assign ecchmatrix[7][220] = 0;
   assign ecchmatrix[8][220] = 1;
   assign ecchmatrix[9][220] = 1;
   assign ecchmatrix[0][221] = 1;
   assign ecchmatrix[1][221] = 0;
   assign ecchmatrix[2][221] = 0;
   assign ecchmatrix[3][221] = 1;
   assign ecchmatrix[4][221] = 0;
   assign ecchmatrix[5][221] = 1;
   assign ecchmatrix[6][221] = 1;
   assign ecchmatrix[7][221] = 1;
   assign ecchmatrix[8][221] = 0;
   assign ecchmatrix[9][221] = 0;
   assign ecchmatrix[0][222] = 1;
   assign ecchmatrix[1][222] = 0;
   assign ecchmatrix[2][222] = 0;
   assign ecchmatrix[3][222] = 1;
   assign ecchmatrix[4][222] = 0;
   assign ecchmatrix[5][222] = 1;
   assign ecchmatrix[6][222] = 1;
   assign ecchmatrix[7][222] = 0;
   assign ecchmatrix[8][222] = 1;
   assign ecchmatrix[9][222] = 0;
   assign ecchmatrix[0][223] = 1;
   assign ecchmatrix[1][223] = 0;
   assign ecchmatrix[2][223] = 0;
   assign ecchmatrix[3][223] = 1;
   assign ecchmatrix[4][223] = 0;
   assign ecchmatrix[5][223] = 1;
   assign ecchmatrix[6][223] = 1;
   assign ecchmatrix[7][223] = 0;
   assign ecchmatrix[8][223] = 0;
   assign ecchmatrix[9][223] = 1;
   assign ecchmatrix[0][224] = 1;
   assign ecchmatrix[1][224] = 0;
   assign ecchmatrix[2][224] = 0;
   assign ecchmatrix[3][224] = 1;
   assign ecchmatrix[4][224] = 0;
   assign ecchmatrix[5][224] = 1;
   assign ecchmatrix[6][224] = 0;
   assign ecchmatrix[7][224] = 1;
   assign ecchmatrix[8][224] = 1;
   assign ecchmatrix[9][224] = 0;
   assign ecchmatrix[0][225] = 1;
   assign ecchmatrix[1][225] = 0;
   assign ecchmatrix[2][225] = 0;
   assign ecchmatrix[3][225] = 1;
   assign ecchmatrix[4][225] = 0;
   assign ecchmatrix[5][225] = 1;
   assign ecchmatrix[6][225] = 0;
   assign ecchmatrix[7][225] = 1;
   assign ecchmatrix[8][225] = 0;
   assign ecchmatrix[9][225] = 1;
   assign ecchmatrix[0][226] = 1;
   assign ecchmatrix[1][226] = 0;
   assign ecchmatrix[2][226] = 0;
   assign ecchmatrix[3][226] = 1;
   assign ecchmatrix[4][226] = 0;
   assign ecchmatrix[5][226] = 1;
   assign ecchmatrix[6][226] = 0;
   assign ecchmatrix[7][226] = 0;
   assign ecchmatrix[8][226] = 1;
   assign ecchmatrix[9][226] = 1;
   assign ecchmatrix[0][227] = 1;
   assign ecchmatrix[1][227] = 0;
   assign ecchmatrix[2][227] = 0;
   assign ecchmatrix[3][227] = 1;
   assign ecchmatrix[4][227] = 0;
   assign ecchmatrix[5][227] = 0;
   assign ecchmatrix[6][227] = 1;
   assign ecchmatrix[7][227] = 1;
   assign ecchmatrix[8][227] = 1;
   assign ecchmatrix[9][227] = 0;
   assign ecchmatrix[0][228] = 1;
   assign ecchmatrix[1][228] = 0;
   assign ecchmatrix[2][228] = 0;
   assign ecchmatrix[3][228] = 1;
   assign ecchmatrix[4][228] = 0;
   assign ecchmatrix[5][228] = 0;
   assign ecchmatrix[6][228] = 1;
   assign ecchmatrix[7][228] = 1;
   assign ecchmatrix[8][228] = 0;
   assign ecchmatrix[9][228] = 1;
   assign ecchmatrix[0][229] = 1;
   assign ecchmatrix[1][229] = 0;
   assign ecchmatrix[2][229] = 0;
   assign ecchmatrix[3][229] = 1;
   assign ecchmatrix[4][229] = 0;
   assign ecchmatrix[5][229] = 0;
   assign ecchmatrix[6][229] = 1;
   assign ecchmatrix[7][229] = 0;
   assign ecchmatrix[8][229] = 1;
   assign ecchmatrix[9][229] = 1;
   assign ecchmatrix[0][230] = 1;
   assign ecchmatrix[1][230] = 0;
   assign ecchmatrix[2][230] = 0;
   assign ecchmatrix[3][230] = 1;
   assign ecchmatrix[4][230] = 0;
   assign ecchmatrix[5][230] = 0;
   assign ecchmatrix[6][230] = 0;
   assign ecchmatrix[7][230] = 1;
   assign ecchmatrix[8][230] = 1;
   assign ecchmatrix[9][230] = 1;
   assign ecchmatrix[0][231] = 1;
   assign ecchmatrix[1][231] = 0;
   assign ecchmatrix[2][231] = 0;
   assign ecchmatrix[3][231] = 0;
   assign ecchmatrix[4][231] = 1;
   assign ecchmatrix[5][231] = 1;
   assign ecchmatrix[6][231] = 1;
   assign ecchmatrix[7][231] = 1;
   assign ecchmatrix[8][231] = 0;
   assign ecchmatrix[9][231] = 0;
   assign ecchmatrix[0][232] = 1;
   assign ecchmatrix[1][232] = 0;
   assign ecchmatrix[2][232] = 0;
   assign ecchmatrix[3][232] = 0;
   assign ecchmatrix[4][232] = 1;
   assign ecchmatrix[5][232] = 1;
   assign ecchmatrix[6][232] = 1;
   assign ecchmatrix[7][232] = 0;
   assign ecchmatrix[8][232] = 1;
   assign ecchmatrix[9][232] = 0;
   assign ecchmatrix[0][233] = 1;
   assign ecchmatrix[1][233] = 0;
   assign ecchmatrix[2][233] = 0;
   assign ecchmatrix[3][233] = 0;
   assign ecchmatrix[4][233] = 1;
   assign ecchmatrix[5][233] = 1;
   assign ecchmatrix[6][233] = 1;
   assign ecchmatrix[7][233] = 0;
   assign ecchmatrix[8][233] = 0;
   assign ecchmatrix[9][233] = 1;
   assign ecchmatrix[0][234] = 1;
   assign ecchmatrix[1][234] = 0;
   assign ecchmatrix[2][234] = 0;
   assign ecchmatrix[3][234] = 0;
   assign ecchmatrix[4][234] = 1;
   assign ecchmatrix[5][234] = 1;
   assign ecchmatrix[6][234] = 0;
   assign ecchmatrix[7][234] = 1;
   assign ecchmatrix[8][234] = 1;
   assign ecchmatrix[9][234] = 0;
   assign ecchmatrix[0][235] = 1;
   assign ecchmatrix[1][235] = 0;
   assign ecchmatrix[2][235] = 0;
   assign ecchmatrix[3][235] = 0;
   assign ecchmatrix[4][235] = 1;
   assign ecchmatrix[5][235] = 1;
   assign ecchmatrix[6][235] = 0;
   assign ecchmatrix[7][235] = 1;
   assign ecchmatrix[8][235] = 0;
   assign ecchmatrix[9][235] = 1;
   assign ecchmatrix[0][236] = 1;
   assign ecchmatrix[1][236] = 0;
   assign ecchmatrix[2][236] = 0;
   assign ecchmatrix[3][236] = 0;
   assign ecchmatrix[4][236] = 1;
   assign ecchmatrix[5][236] = 1;
   assign ecchmatrix[6][236] = 0;
   assign ecchmatrix[7][236] = 0;
   assign ecchmatrix[8][236] = 1;
   assign ecchmatrix[9][236] = 1;
   assign ecchmatrix[0][237] = 1;
   assign ecchmatrix[1][237] = 0;
   assign ecchmatrix[2][237] = 0;
   assign ecchmatrix[3][237] = 0;
   assign ecchmatrix[4][237] = 1;
   assign ecchmatrix[5][237] = 0;
   assign ecchmatrix[6][237] = 1;
   assign ecchmatrix[7][237] = 1;
   assign ecchmatrix[8][237] = 1;
   assign ecchmatrix[9][237] = 0;
   assign ecchmatrix[0][238] = 1;
   assign ecchmatrix[1][238] = 0;
   assign ecchmatrix[2][238] = 0;
   assign ecchmatrix[3][238] = 0;
   assign ecchmatrix[4][238] = 1;
   assign ecchmatrix[5][238] = 0;
   assign ecchmatrix[6][238] = 1;
   assign ecchmatrix[7][238] = 1;
   assign ecchmatrix[8][238] = 0;
   assign ecchmatrix[9][238] = 1;
   assign ecchmatrix[0][239] = 1;
   assign ecchmatrix[1][239] = 0;
   assign ecchmatrix[2][239] = 0;
   assign ecchmatrix[3][239] = 0;
   assign ecchmatrix[4][239] = 1;
   assign ecchmatrix[5][239] = 0;
   assign ecchmatrix[6][239] = 1;
   assign ecchmatrix[7][239] = 0;
   assign ecchmatrix[8][239] = 1;
   assign ecchmatrix[9][239] = 1;
   assign ecchmatrix[0][240] = 1;
   assign ecchmatrix[1][240] = 0;
   assign ecchmatrix[2][240] = 0;
   assign ecchmatrix[3][240] = 0;
   assign ecchmatrix[4][240] = 1;
   assign ecchmatrix[5][240] = 0;
   assign ecchmatrix[6][240] = 0;
   assign ecchmatrix[7][240] = 1;
   assign ecchmatrix[8][240] = 1;
   assign ecchmatrix[9][240] = 1;
   assign ecchmatrix[0][241] = 1;
   assign ecchmatrix[1][241] = 0;
   assign ecchmatrix[2][241] = 0;
   assign ecchmatrix[3][241] = 0;
   assign ecchmatrix[4][241] = 0;
   assign ecchmatrix[5][241] = 1;
   assign ecchmatrix[6][241] = 1;
   assign ecchmatrix[7][241] = 1;
   assign ecchmatrix[8][241] = 1;
   assign ecchmatrix[9][241] = 0;
   assign ecchmatrix[0][242] = 1;
   assign ecchmatrix[1][242] = 0;
   assign ecchmatrix[2][242] = 0;
   assign ecchmatrix[3][242] = 0;
   assign ecchmatrix[4][242] = 0;
   assign ecchmatrix[5][242] = 1;
   assign ecchmatrix[6][242] = 1;
   assign ecchmatrix[7][242] = 1;
   assign ecchmatrix[8][242] = 0;
   assign ecchmatrix[9][242] = 1;
   assign ecchmatrix[0][243] = 1;
   assign ecchmatrix[1][243] = 0;
   assign ecchmatrix[2][243] = 0;
   assign ecchmatrix[3][243] = 0;
   assign ecchmatrix[4][243] = 0;
   assign ecchmatrix[5][243] = 1;
   assign ecchmatrix[6][243] = 1;
   assign ecchmatrix[7][243] = 0;
   assign ecchmatrix[8][243] = 1;
   assign ecchmatrix[9][243] = 1;
   assign ecchmatrix[0][244] = 1;
   assign ecchmatrix[1][244] = 0;
   assign ecchmatrix[2][244] = 0;
   assign ecchmatrix[3][244] = 0;
   assign ecchmatrix[4][244] = 0;
   assign ecchmatrix[5][244] = 1;
   assign ecchmatrix[6][244] = 0;
   assign ecchmatrix[7][244] = 1;
   assign ecchmatrix[8][244] = 1;
   assign ecchmatrix[9][244] = 1;
   assign ecchmatrix[0][245] = 1;
   assign ecchmatrix[1][245] = 0;
   assign ecchmatrix[2][245] = 0;
   assign ecchmatrix[3][245] = 0;
   assign ecchmatrix[4][245] = 0;
   assign ecchmatrix[5][245] = 0;
   assign ecchmatrix[6][245] = 1;
   assign ecchmatrix[7][245] = 1;
   assign ecchmatrix[8][245] = 1;
   assign ecchmatrix[9][245] = 1;
   assign ecchmatrix[0][246] = 0;
   assign ecchmatrix[1][246] = 1;
   assign ecchmatrix[2][246] = 1;
   assign ecchmatrix[3][246] = 1;
   assign ecchmatrix[4][246] = 1;
   assign ecchmatrix[5][246] = 1;
   assign ecchmatrix[6][246] = 0;
   assign ecchmatrix[7][246] = 0;
   assign ecchmatrix[8][246] = 0;
   assign ecchmatrix[9][246] = 0;
   assign ecchmatrix[0][247] = 0;
   assign ecchmatrix[1][247] = 1;
   assign ecchmatrix[2][247] = 1;
   assign ecchmatrix[3][247] = 1;
   assign ecchmatrix[4][247] = 1;
   assign ecchmatrix[5][247] = 0;
   assign ecchmatrix[6][247] = 1;
   assign ecchmatrix[7][247] = 0;
   assign ecchmatrix[8][247] = 0;
   assign ecchmatrix[9][247] = 0;
   assign ecchmatrix[0][248] = 0;
   assign ecchmatrix[1][248] = 1;
   assign ecchmatrix[2][248] = 1;
   assign ecchmatrix[3][248] = 1;
   assign ecchmatrix[4][248] = 1;
   assign ecchmatrix[5][248] = 0;
   assign ecchmatrix[6][248] = 0;
   assign ecchmatrix[7][248] = 1;
   assign ecchmatrix[8][248] = 0;
   assign ecchmatrix[9][248] = 0;
   assign ecchmatrix[0][249] = 0;
   assign ecchmatrix[1][249] = 1;
   assign ecchmatrix[2][249] = 1;
   assign ecchmatrix[3][249] = 1;
   assign ecchmatrix[4][249] = 1;
   assign ecchmatrix[5][249] = 0;
   assign ecchmatrix[6][249] = 0;
   assign ecchmatrix[7][249] = 0;
   assign ecchmatrix[8][249] = 1;
   assign ecchmatrix[9][249] = 0;
   assign ecchmatrix[0][250] = 0;
   assign ecchmatrix[1][250] = 1;
   assign ecchmatrix[2][250] = 1;
   assign ecchmatrix[3][250] = 1;
   assign ecchmatrix[4][250] = 1;
   assign ecchmatrix[5][250] = 0;
   assign ecchmatrix[6][250] = 0;
   assign ecchmatrix[7][250] = 0;
   assign ecchmatrix[8][250] = 0;
   assign ecchmatrix[9][250] = 1;
   assign ecchmatrix[0][251] = 0;
   assign ecchmatrix[1][251] = 1;
   assign ecchmatrix[2][251] = 1;
   assign ecchmatrix[3][251] = 1;
   assign ecchmatrix[4][251] = 0;
   assign ecchmatrix[5][251] = 1;
   assign ecchmatrix[6][251] = 1;
   assign ecchmatrix[7][251] = 0;
   assign ecchmatrix[8][251] = 0;
   assign ecchmatrix[9][251] = 0;
   assign ecchmatrix[0][252] = 0;
   assign ecchmatrix[1][252] = 1;
   assign ecchmatrix[2][252] = 1;
   assign ecchmatrix[3][252] = 1;
   assign ecchmatrix[4][252] = 0;
   assign ecchmatrix[5][252] = 1;
   assign ecchmatrix[6][252] = 0;
   assign ecchmatrix[7][252] = 1;
   assign ecchmatrix[8][252] = 0;
   assign ecchmatrix[9][252] = 0;
   assign ecchmatrix[0][253] = 0;
   assign ecchmatrix[1][253] = 1;
   assign ecchmatrix[2][253] = 1;
   assign ecchmatrix[3][253] = 1;
   assign ecchmatrix[4][253] = 0;
   assign ecchmatrix[5][253] = 1;
   assign ecchmatrix[6][253] = 0;
   assign ecchmatrix[7][253] = 0;
   assign ecchmatrix[8][253] = 1;
   assign ecchmatrix[9][253] = 0;
   assign ecchmatrix[0][254] = 0;
   assign ecchmatrix[1][254] = 1;
   assign ecchmatrix[2][254] = 1;
   assign ecchmatrix[3][254] = 1;
   assign ecchmatrix[4][254] = 0;
   assign ecchmatrix[5][254] = 1;
   assign ecchmatrix[6][254] = 0;
   assign ecchmatrix[7][254] = 0;
   assign ecchmatrix[8][254] = 0;
   assign ecchmatrix[9][254] = 1;
   assign ecchmatrix[0][255] = 0;
   assign ecchmatrix[1][255] = 1;
   assign ecchmatrix[2][255] = 1;
   assign ecchmatrix[3][255] = 1;
   assign ecchmatrix[4][255] = 0;
   assign ecchmatrix[5][255] = 0;
   assign ecchmatrix[6][255] = 1;
   assign ecchmatrix[7][255] = 1;
   assign ecchmatrix[8][255] = 0;
   assign ecchmatrix[9][255] = 0;
   assign ecchmatrix[0][256] = 0;
   assign ecchmatrix[1][256] = 1;
   assign ecchmatrix[2][256] = 1;
   assign ecchmatrix[3][256] = 1;
   assign ecchmatrix[4][256] = 0;
   assign ecchmatrix[5][256] = 0;
   assign ecchmatrix[6][256] = 1;
   assign ecchmatrix[7][256] = 0;
   assign ecchmatrix[8][256] = 1;
   assign ecchmatrix[9][256] = 0;
   assign ecchmatrix[0][257] = 0;
   assign ecchmatrix[1][257] = 1;
   assign ecchmatrix[2][257] = 1;
   assign ecchmatrix[3][257] = 1;
   assign ecchmatrix[4][257] = 0;
   assign ecchmatrix[5][257] = 0;
   assign ecchmatrix[6][257] = 1;
   assign ecchmatrix[7][257] = 0;
   assign ecchmatrix[8][257] = 0;
   assign ecchmatrix[9][257] = 1;
   assign ecchmatrix[0][258] = 0;
   assign ecchmatrix[1][258] = 1;
   assign ecchmatrix[2][258] = 1;
   assign ecchmatrix[3][258] = 1;
   assign ecchmatrix[4][258] = 0;
   assign ecchmatrix[5][258] = 0;
   assign ecchmatrix[6][258] = 0;
   assign ecchmatrix[7][258] = 1;
   assign ecchmatrix[8][258] = 1;
   assign ecchmatrix[9][258] = 0;
   assign ecchmatrix[0][259] = 0;
   assign ecchmatrix[1][259] = 1;
   assign ecchmatrix[2][259] = 1;
   assign ecchmatrix[3][259] = 1;
   assign ecchmatrix[4][259] = 0;
   assign ecchmatrix[5][259] = 0;
   assign ecchmatrix[6][259] = 0;
   assign ecchmatrix[7][259] = 1;
   assign ecchmatrix[8][259] = 0;
   assign ecchmatrix[9][259] = 1;
   assign ecchmatrix[0][260] = 0;
   assign ecchmatrix[1][260] = 1;
   assign ecchmatrix[2][260] = 1;
   assign ecchmatrix[3][260] = 1;
   assign ecchmatrix[4][260] = 0;
   assign ecchmatrix[5][260] = 0;
   assign ecchmatrix[6][260] = 0;
   assign ecchmatrix[7][260] = 0;
   assign ecchmatrix[8][260] = 1;
   assign ecchmatrix[9][260] = 1;
   assign ecchmatrix[0][261] = 0;
   assign ecchmatrix[1][261] = 1;
   assign ecchmatrix[2][261] = 1;
   assign ecchmatrix[3][261] = 0;
   assign ecchmatrix[4][261] = 1;
   assign ecchmatrix[5][261] = 1;
   assign ecchmatrix[6][261] = 1;
   assign ecchmatrix[7][261] = 0;
   assign ecchmatrix[8][261] = 0;
   assign ecchmatrix[9][261] = 0;
   assign ecchmatrix[0][262] = 0;
   assign ecchmatrix[1][262] = 1;
   assign ecchmatrix[2][262] = 1;
   assign ecchmatrix[3][262] = 0;
   assign ecchmatrix[4][262] = 1;
   assign ecchmatrix[5][262] = 1;
   assign ecchmatrix[6][262] = 0;
   assign ecchmatrix[7][262] = 1;
   assign ecchmatrix[8][262] = 0;
   assign ecchmatrix[9][262] = 0;
   assign ecchmatrix[0][263] = 0;
   assign ecchmatrix[1][263] = 1;
   assign ecchmatrix[2][263] = 1;
   assign ecchmatrix[3][263] = 0;
   assign ecchmatrix[4][263] = 1;
   assign ecchmatrix[5][263] = 1;
   assign ecchmatrix[6][263] = 0;
   assign ecchmatrix[7][263] = 0;
   assign ecchmatrix[8][263] = 1;
   assign ecchmatrix[9][263] = 0;
   assign ecchmatrix[0][264] = 0;
   assign ecchmatrix[1][264] = 1;
   assign ecchmatrix[2][264] = 1;
   assign ecchmatrix[3][264] = 0;
   assign ecchmatrix[4][264] = 1;
   assign ecchmatrix[5][264] = 1;
   assign ecchmatrix[6][264] = 0;
   assign ecchmatrix[7][264] = 0;
   assign ecchmatrix[8][264] = 0;
   assign ecchmatrix[9][264] = 1;
   assign ecchmatrix[0][265] = 0;
   assign ecchmatrix[1][265] = 1;
   assign ecchmatrix[2][265] = 1;
   assign ecchmatrix[3][265] = 0;
   assign ecchmatrix[4][265] = 1;
   assign ecchmatrix[5][265] = 0;
   assign ecchmatrix[6][265] = 1;
   assign ecchmatrix[7][265] = 1;
   assign ecchmatrix[8][265] = 0;
   assign ecchmatrix[9][265] = 0;
   assign ecchmatrix[0][266] = 0;
   assign ecchmatrix[1][266] = 1;
   assign ecchmatrix[2][266] = 1;
   assign ecchmatrix[3][266] = 0;
   assign ecchmatrix[4][266] = 1;
   assign ecchmatrix[5][266] = 0;
   assign ecchmatrix[6][266] = 1;
   assign ecchmatrix[7][266] = 0;
   assign ecchmatrix[8][266] = 1;
   assign ecchmatrix[9][266] = 0;
   assign ecchmatrix[0][267] = 0;
   assign ecchmatrix[1][267] = 1;
   assign ecchmatrix[2][267] = 1;
   assign ecchmatrix[3][267] = 0;
   assign ecchmatrix[4][267] = 1;
   assign ecchmatrix[5][267] = 0;
   assign ecchmatrix[6][267] = 1;
   assign ecchmatrix[7][267] = 0;
   assign ecchmatrix[8][267] = 0;
   assign ecchmatrix[9][267] = 1;
   assign ecchmatrix[0][268] = 0;
   assign ecchmatrix[1][268] = 1;
   assign ecchmatrix[2][268] = 1;
   assign ecchmatrix[3][268] = 0;
   assign ecchmatrix[4][268] = 1;
   assign ecchmatrix[5][268] = 0;
   assign ecchmatrix[6][268] = 0;
   assign ecchmatrix[7][268] = 1;
   assign ecchmatrix[8][268] = 1;
   assign ecchmatrix[9][268] = 0;
   assign ecchmatrix[0][269] = 0;
   assign ecchmatrix[1][269] = 1;
   assign ecchmatrix[2][269] = 1;
   assign ecchmatrix[3][269] = 0;
   assign ecchmatrix[4][269] = 1;
   assign ecchmatrix[5][269] = 0;
   assign ecchmatrix[6][269] = 0;
   assign ecchmatrix[7][269] = 1;
   assign ecchmatrix[8][269] = 0;
   assign ecchmatrix[9][269] = 1;
   assign ecchmatrix[0][270] = 0;
   assign ecchmatrix[1][270] = 1;
   assign ecchmatrix[2][270] = 1;
   assign ecchmatrix[3][270] = 0;
   assign ecchmatrix[4][270] = 1;
   assign ecchmatrix[5][270] = 0;
   assign ecchmatrix[6][270] = 0;
   assign ecchmatrix[7][270] = 0;
   assign ecchmatrix[8][270] = 1;
   assign ecchmatrix[9][270] = 1;
   assign ecchmatrix[0][271] = 0;
   assign ecchmatrix[1][271] = 1;
   assign ecchmatrix[2][271] = 1;
   assign ecchmatrix[3][271] = 0;
   assign ecchmatrix[4][271] = 0;
   assign ecchmatrix[5][271] = 1;
   assign ecchmatrix[6][271] = 1;
   assign ecchmatrix[7][271] = 1;
   assign ecchmatrix[8][271] = 0;
   assign ecchmatrix[9][271] = 0;
   assign ecchmatrix[0][272] = 0;
   assign ecchmatrix[1][272] = 1;
   assign ecchmatrix[2][272] = 1;
   assign ecchmatrix[3][272] = 0;
   assign ecchmatrix[4][272] = 0;
   assign ecchmatrix[5][272] = 1;
   assign ecchmatrix[6][272] = 1;
   assign ecchmatrix[7][272] = 0;
   assign ecchmatrix[8][272] = 1;
   assign ecchmatrix[9][272] = 0;
   assign ecchmatrix[0][273] = 0;
   assign ecchmatrix[1][273] = 1;
   assign ecchmatrix[2][273] = 1;
   assign ecchmatrix[3][273] = 0;
   assign ecchmatrix[4][273] = 0;
   assign ecchmatrix[5][273] = 1;
   assign ecchmatrix[6][273] = 1;
   assign ecchmatrix[7][273] = 0;
   assign ecchmatrix[8][273] = 0;
   assign ecchmatrix[9][273] = 1;
   assign ecchmatrix[0][274] = 0;
   assign ecchmatrix[1][274] = 1;
   assign ecchmatrix[2][274] = 1;
   assign ecchmatrix[3][274] = 0;
   assign ecchmatrix[4][274] = 0;
   assign ecchmatrix[5][274] = 1;
   assign ecchmatrix[6][274] = 0;
   assign ecchmatrix[7][274] = 1;
   assign ecchmatrix[8][274] = 1;
   assign ecchmatrix[9][274] = 0;
   assign ecchmatrix[0][275] = 0;
   assign ecchmatrix[1][275] = 1;
   assign ecchmatrix[2][275] = 1;
   assign ecchmatrix[3][275] = 0;
   assign ecchmatrix[4][275] = 0;
   assign ecchmatrix[5][275] = 1;
   assign ecchmatrix[6][275] = 0;
   assign ecchmatrix[7][275] = 1;
   assign ecchmatrix[8][275] = 0;
   assign ecchmatrix[9][275] = 1;
   assign ecchmatrix[0][276] = 0;
   assign ecchmatrix[1][276] = 1;
   assign ecchmatrix[2][276] = 1;
   assign ecchmatrix[3][276] = 0;
   assign ecchmatrix[4][276] = 0;
   assign ecchmatrix[5][276] = 1;
   assign ecchmatrix[6][276] = 0;
   assign ecchmatrix[7][276] = 0;
   assign ecchmatrix[8][276] = 1;
   assign ecchmatrix[9][276] = 1;
   assign ecchmatrix[0][277] = 0;
   assign ecchmatrix[1][277] = 1;
   assign ecchmatrix[2][277] = 1;
   assign ecchmatrix[3][277] = 0;
   assign ecchmatrix[4][277] = 0;
   assign ecchmatrix[5][277] = 0;
   assign ecchmatrix[6][277] = 1;
   assign ecchmatrix[7][277] = 1;
   assign ecchmatrix[8][277] = 1;
   assign ecchmatrix[9][277] = 0;
   assign ecchmatrix[0][278] = 0;
   assign ecchmatrix[1][278] = 1;
   assign ecchmatrix[2][278] = 1;
   assign ecchmatrix[3][278] = 0;
   assign ecchmatrix[4][278] = 0;
   assign ecchmatrix[5][278] = 0;
   assign ecchmatrix[6][278] = 1;
   assign ecchmatrix[7][278] = 1;
   assign ecchmatrix[8][278] = 0;
   assign ecchmatrix[9][278] = 1;
   assign ecchmatrix[0][279] = 0;
   assign ecchmatrix[1][279] = 1;
   assign ecchmatrix[2][279] = 1;
   assign ecchmatrix[3][279] = 0;
   assign ecchmatrix[4][279] = 0;
   assign ecchmatrix[5][279] = 0;
   assign ecchmatrix[6][279] = 1;
   assign ecchmatrix[7][279] = 0;
   assign ecchmatrix[8][279] = 1;
   assign ecchmatrix[9][279] = 1;
   assign ecchmatrix[0][280] = 0;
   assign ecchmatrix[1][280] = 1;
   assign ecchmatrix[2][280] = 1;
   assign ecchmatrix[3][280] = 0;
   assign ecchmatrix[4][280] = 0;
   assign ecchmatrix[5][280] = 0;
   assign ecchmatrix[6][280] = 0;
   assign ecchmatrix[7][280] = 1;
   assign ecchmatrix[8][280] = 1;
   assign ecchmatrix[9][280] = 1;
   assign ecchmatrix[0][281] = 0;
   assign ecchmatrix[1][281] = 1;
   assign ecchmatrix[2][281] = 0;
   assign ecchmatrix[3][281] = 1;
   assign ecchmatrix[4][281] = 1;
   assign ecchmatrix[5][281] = 1;
   assign ecchmatrix[6][281] = 1;
   assign ecchmatrix[7][281] = 0;
   assign ecchmatrix[8][281] = 0;
   assign ecchmatrix[9][281] = 0;
   assign ecchmatrix[0][282] = 0;
   assign ecchmatrix[1][282] = 1;
   assign ecchmatrix[2][282] = 0;
   assign ecchmatrix[3][282] = 1;
   assign ecchmatrix[4][282] = 1;
   assign ecchmatrix[5][282] = 1;
   assign ecchmatrix[6][282] = 0;
   assign ecchmatrix[7][282] = 1;
   assign ecchmatrix[8][282] = 0;
   assign ecchmatrix[9][282] = 0;
   assign ecchmatrix[0][283] = 0;
   assign ecchmatrix[1][283] = 1;
   assign ecchmatrix[2][283] = 0;
   assign ecchmatrix[3][283] = 1;
   assign ecchmatrix[4][283] = 1;
   assign ecchmatrix[5][283] = 1;
   assign ecchmatrix[6][283] = 0;
   assign ecchmatrix[7][283] = 0;
   assign ecchmatrix[8][283] = 1;
   assign ecchmatrix[9][283] = 0;
   assign ecchmatrix[0][284] = 0;
   assign ecchmatrix[1][284] = 1;
   assign ecchmatrix[2][284] = 0;
   assign ecchmatrix[3][284] = 1;
   assign ecchmatrix[4][284] = 1;
   assign ecchmatrix[5][284] = 1;
   assign ecchmatrix[6][284] = 0;
   assign ecchmatrix[7][284] = 0;
   assign ecchmatrix[8][284] = 0;
   assign ecchmatrix[9][284] = 1;
   assign ecchmatrix[0][285] = 0;
   assign ecchmatrix[1][285] = 1;
   assign ecchmatrix[2][285] = 0;
   assign ecchmatrix[3][285] = 1;
   assign ecchmatrix[4][285] = 1;
   assign ecchmatrix[5][285] = 0;
   assign ecchmatrix[6][285] = 1;
   assign ecchmatrix[7][285] = 1;
   assign ecchmatrix[8][285] = 0;
   assign ecchmatrix[9][285] = 0;
   assign ecchmatrix[0][286] = 0;
   assign ecchmatrix[1][286] = 1;
   assign ecchmatrix[2][286] = 0;
   assign ecchmatrix[3][286] = 1;
   assign ecchmatrix[4][286] = 1;
   assign ecchmatrix[5][286] = 0;
   assign ecchmatrix[6][286] = 1;
   assign ecchmatrix[7][286] = 0;
   assign ecchmatrix[8][286] = 1;
   assign ecchmatrix[9][286] = 0;
   assign ecchmatrix[0][287] = 0;
   assign ecchmatrix[1][287] = 1;
   assign ecchmatrix[2][287] = 0;
   assign ecchmatrix[3][287] = 1;
   assign ecchmatrix[4][287] = 1;
   assign ecchmatrix[5][287] = 0;
   assign ecchmatrix[6][287] = 1;
   assign ecchmatrix[7][287] = 0;
   assign ecchmatrix[8][287] = 0;
   assign ecchmatrix[9][287] = 1;
   assign ecchmatrix[0][288] = 0;
   assign ecchmatrix[1][288] = 1;
   assign ecchmatrix[2][288] = 0;
   assign ecchmatrix[3][288] = 1;
   assign ecchmatrix[4][288] = 1;
   assign ecchmatrix[5][288] = 0;
   assign ecchmatrix[6][288] = 0;
   assign ecchmatrix[7][288] = 1;
   assign ecchmatrix[8][288] = 1;
   assign ecchmatrix[9][288] = 0;
   assign ecchmatrix[0][289] = 0;
   assign ecchmatrix[1][289] = 1;
   assign ecchmatrix[2][289] = 0;
   assign ecchmatrix[3][289] = 1;
   assign ecchmatrix[4][289] = 1;
   assign ecchmatrix[5][289] = 0;
   assign ecchmatrix[6][289] = 0;
   assign ecchmatrix[7][289] = 1;
   assign ecchmatrix[8][289] = 0;
   assign ecchmatrix[9][289] = 1;
   assign ecchmatrix[0][290] = 0;
   assign ecchmatrix[1][290] = 1;
   assign ecchmatrix[2][290] = 0;
   assign ecchmatrix[3][290] = 1;
   assign ecchmatrix[4][290] = 1;
   assign ecchmatrix[5][290] = 0;
   assign ecchmatrix[6][290] = 0;
   assign ecchmatrix[7][290] = 0;
   assign ecchmatrix[8][290] = 1;
   assign ecchmatrix[9][290] = 1;
   assign ecchmatrix[0][291] = 0;
   assign ecchmatrix[1][291] = 1;
   assign ecchmatrix[2][291] = 0;
   assign ecchmatrix[3][291] = 1;
   assign ecchmatrix[4][291] = 0;
   assign ecchmatrix[5][291] = 1;
   assign ecchmatrix[6][291] = 1;
   assign ecchmatrix[7][291] = 1;
   assign ecchmatrix[8][291] = 0;
   assign ecchmatrix[9][291] = 0;
   assign ecchmatrix[0][292] = 0;
   assign ecchmatrix[1][292] = 1;
   assign ecchmatrix[2][292] = 0;
   assign ecchmatrix[3][292] = 1;
   assign ecchmatrix[4][292] = 0;
   assign ecchmatrix[5][292] = 1;
   assign ecchmatrix[6][292] = 1;
   assign ecchmatrix[7][292] = 0;
   assign ecchmatrix[8][292] = 1;
   assign ecchmatrix[9][292] = 0;
   assign ecchmatrix[0][293] = 0;
   assign ecchmatrix[1][293] = 1;
   assign ecchmatrix[2][293] = 0;
   assign ecchmatrix[3][293] = 1;
   assign ecchmatrix[4][293] = 0;
   assign ecchmatrix[5][293] = 1;
   assign ecchmatrix[6][293] = 1;
   assign ecchmatrix[7][293] = 0;
   assign ecchmatrix[8][293] = 0;
   assign ecchmatrix[9][293] = 1;
   assign ecchmatrix[0][294] = 0;
   assign ecchmatrix[1][294] = 1;
   assign ecchmatrix[2][294] = 0;
   assign ecchmatrix[3][294] = 1;
   assign ecchmatrix[4][294] = 0;
   assign ecchmatrix[5][294] = 1;
   assign ecchmatrix[6][294] = 0;
   assign ecchmatrix[7][294] = 1;
   assign ecchmatrix[8][294] = 1;
   assign ecchmatrix[9][294] = 0;
   assign ecchmatrix[0][295] = 0;
   assign ecchmatrix[1][295] = 1;
   assign ecchmatrix[2][295] = 0;
   assign ecchmatrix[3][295] = 1;
   assign ecchmatrix[4][295] = 0;
   assign ecchmatrix[5][295] = 1;
   assign ecchmatrix[6][295] = 0;
   assign ecchmatrix[7][295] = 1;
   assign ecchmatrix[8][295] = 0;
   assign ecchmatrix[9][295] = 1;
   assign ecchmatrix[0][296] = 0;
   assign ecchmatrix[1][296] = 1;
   assign ecchmatrix[2][296] = 0;
   assign ecchmatrix[3][296] = 1;
   assign ecchmatrix[4][296] = 0;
   assign ecchmatrix[5][296] = 1;
   assign ecchmatrix[6][296] = 0;
   assign ecchmatrix[7][296] = 0;
   assign ecchmatrix[8][296] = 1;
   assign ecchmatrix[9][296] = 1;
   assign ecchmatrix[0][297] = 0;
   assign ecchmatrix[1][297] = 1;
   assign ecchmatrix[2][297] = 0;
   assign ecchmatrix[3][297] = 1;
   assign ecchmatrix[4][297] = 0;
   assign ecchmatrix[5][297] = 0;
   assign ecchmatrix[6][297] = 1;
   assign ecchmatrix[7][297] = 1;
   assign ecchmatrix[8][297] = 1;
   assign ecchmatrix[9][297] = 0;
   assign ecchmatrix[0][298] = 0;
   assign ecchmatrix[1][298] = 1;
   assign ecchmatrix[2][298] = 0;
   assign ecchmatrix[3][298] = 1;
   assign ecchmatrix[4][298] = 0;
   assign ecchmatrix[5][298] = 0;
   assign ecchmatrix[6][298] = 1;
   assign ecchmatrix[7][298] = 1;
   assign ecchmatrix[8][298] = 0;
   assign ecchmatrix[9][298] = 1;
   assign ecchmatrix[0][299] = 0;
   assign ecchmatrix[1][299] = 1;
   assign ecchmatrix[2][299] = 0;
   assign ecchmatrix[3][299] = 1;
   assign ecchmatrix[4][299] = 0;
   assign ecchmatrix[5][299] = 0;
   assign ecchmatrix[6][299] = 1;
   assign ecchmatrix[7][299] = 0;
   assign ecchmatrix[8][299] = 1;
   assign ecchmatrix[9][299] = 1;
   assign ecchmatrix[0][300] = 0;
   assign ecchmatrix[1][300] = 1;
   assign ecchmatrix[2][300] = 0;
   assign ecchmatrix[3][300] = 1;
   assign ecchmatrix[4][300] = 0;
   assign ecchmatrix[5][300] = 0;
   assign ecchmatrix[6][300] = 0;
   assign ecchmatrix[7][300] = 1;
   assign ecchmatrix[8][300] = 1;
   assign ecchmatrix[9][300] = 1;
   assign ecchmatrix[0][301] = 0;
   assign ecchmatrix[1][301] = 1;
   assign ecchmatrix[2][301] = 0;
   assign ecchmatrix[3][301] = 0;
   assign ecchmatrix[4][301] = 1;
   assign ecchmatrix[5][301] = 1;
   assign ecchmatrix[6][301] = 1;
   assign ecchmatrix[7][301] = 1;
   assign ecchmatrix[8][301] = 0;
   assign ecchmatrix[9][301] = 0;
   assign ecchmatrix[0][302] = 0;
   assign ecchmatrix[1][302] = 1;
   assign ecchmatrix[2][302] = 0;
   assign ecchmatrix[3][302] = 0;
   assign ecchmatrix[4][302] = 1;
   assign ecchmatrix[5][302] = 1;
   assign ecchmatrix[6][302] = 1;
   assign ecchmatrix[7][302] = 0;
   assign ecchmatrix[8][302] = 1;
   assign ecchmatrix[9][302] = 0;
   assign ecchmatrix[0][303] = 0;
   assign ecchmatrix[1][303] = 1;
   assign ecchmatrix[2][303] = 0;
   assign ecchmatrix[3][303] = 0;
   assign ecchmatrix[4][303] = 1;
   assign ecchmatrix[5][303] = 1;
   assign ecchmatrix[6][303] = 1;
   assign ecchmatrix[7][303] = 0;
   assign ecchmatrix[8][303] = 0;
   assign ecchmatrix[9][303] = 1;
   assign ecchmatrix[0][304] = 0;
   assign ecchmatrix[1][304] = 1;
   assign ecchmatrix[2][304] = 0;
   assign ecchmatrix[3][304] = 0;
   assign ecchmatrix[4][304] = 1;
   assign ecchmatrix[5][304] = 1;
   assign ecchmatrix[6][304] = 0;
   assign ecchmatrix[7][304] = 1;
   assign ecchmatrix[8][304] = 1;
   assign ecchmatrix[9][304] = 0;
   assign ecchmatrix[0][305] = 0;
   assign ecchmatrix[1][305] = 1;
   assign ecchmatrix[2][305] = 0;
   assign ecchmatrix[3][305] = 0;
   assign ecchmatrix[4][305] = 1;
   assign ecchmatrix[5][305] = 1;
   assign ecchmatrix[6][305] = 0;
   assign ecchmatrix[7][305] = 1;
   assign ecchmatrix[8][305] = 0;
   assign ecchmatrix[9][305] = 1;
   assign ecchmatrix[0][306] = 0;
   assign ecchmatrix[1][306] = 1;
   assign ecchmatrix[2][306] = 0;
   assign ecchmatrix[3][306] = 0;
   assign ecchmatrix[4][306] = 1;
   assign ecchmatrix[5][306] = 1;
   assign ecchmatrix[6][306] = 0;
   assign ecchmatrix[7][306] = 0;
   assign ecchmatrix[8][306] = 1;
   assign ecchmatrix[9][306] = 1;
   assign ecchmatrix[0][307] = 0;
   assign ecchmatrix[1][307] = 1;
   assign ecchmatrix[2][307] = 0;
   assign ecchmatrix[3][307] = 0;
   assign ecchmatrix[4][307] = 1;
   assign ecchmatrix[5][307] = 0;
   assign ecchmatrix[6][307] = 1;
   assign ecchmatrix[7][307] = 1;
   assign ecchmatrix[8][307] = 1;
   assign ecchmatrix[9][307] = 0;
   assign ecchmatrix[0][308] = 0;
   assign ecchmatrix[1][308] = 1;
   assign ecchmatrix[2][308] = 0;
   assign ecchmatrix[3][308] = 0;
   assign ecchmatrix[4][308] = 1;
   assign ecchmatrix[5][308] = 0;
   assign ecchmatrix[6][308] = 1;
   assign ecchmatrix[7][308] = 1;
   assign ecchmatrix[8][308] = 0;
   assign ecchmatrix[9][308] = 1;
   assign ecchmatrix[0][309] = 0;
   assign ecchmatrix[1][309] = 1;
   assign ecchmatrix[2][309] = 0;
   assign ecchmatrix[3][309] = 0;
   assign ecchmatrix[4][309] = 1;
   assign ecchmatrix[5][309] = 0;
   assign ecchmatrix[6][309] = 1;
   assign ecchmatrix[7][309] = 0;
   assign ecchmatrix[8][309] = 1;
   assign ecchmatrix[9][309] = 1;
   assign ecchmatrix[0][310] = 0;
   assign ecchmatrix[1][310] = 1;
   assign ecchmatrix[2][310] = 0;
   assign ecchmatrix[3][310] = 0;
   assign ecchmatrix[4][310] = 1;
   assign ecchmatrix[5][310] = 0;
   assign ecchmatrix[6][310] = 0;
   assign ecchmatrix[7][310] = 1;
   assign ecchmatrix[8][310] = 1;
   assign ecchmatrix[9][310] = 1;
   assign ecchmatrix[0][311] = 0;
   assign ecchmatrix[1][311] = 1;
   assign ecchmatrix[2][311] = 0;
   assign ecchmatrix[3][311] = 0;
   assign ecchmatrix[4][311] = 0;
   assign ecchmatrix[5][311] = 1;
   assign ecchmatrix[6][311] = 1;
   assign ecchmatrix[7][311] = 1;
   assign ecchmatrix[8][311] = 1;
   assign ecchmatrix[9][311] = 0;
   assign ecchmatrix[0][312] = 0;
   assign ecchmatrix[1][312] = 1;
   assign ecchmatrix[2][312] = 0;
   assign ecchmatrix[3][312] = 0;
   assign ecchmatrix[4][312] = 0;
   assign ecchmatrix[5][312] = 1;
   assign ecchmatrix[6][312] = 1;
   assign ecchmatrix[7][312] = 1;
   assign ecchmatrix[8][312] = 0;
   assign ecchmatrix[9][312] = 1;
   assign ecchmatrix[0][313] = 0;
   assign ecchmatrix[1][313] = 1;
   assign ecchmatrix[2][313] = 0;
   assign ecchmatrix[3][313] = 0;
   assign ecchmatrix[4][313] = 0;
   assign ecchmatrix[5][313] = 1;
   assign ecchmatrix[6][313] = 1;
   assign ecchmatrix[7][313] = 0;
   assign ecchmatrix[8][313] = 1;
   assign ecchmatrix[9][313] = 1;
   assign ecchmatrix[0][314] = 0;
   assign ecchmatrix[1][314] = 1;
   assign ecchmatrix[2][314] = 0;
   assign ecchmatrix[3][314] = 0;
   assign ecchmatrix[4][314] = 0;
   assign ecchmatrix[5][314] = 1;
   assign ecchmatrix[6][314] = 0;
   assign ecchmatrix[7][314] = 1;
   assign ecchmatrix[8][314] = 1;
   assign ecchmatrix[9][314] = 1;
   assign ecchmatrix[0][315] = 0;
   assign ecchmatrix[1][315] = 1;
   assign ecchmatrix[2][315] = 0;
   assign ecchmatrix[3][315] = 0;
   assign ecchmatrix[4][315] = 0;
   assign ecchmatrix[5][315] = 0;
   assign ecchmatrix[6][315] = 1;
   assign ecchmatrix[7][315] = 1;
   assign ecchmatrix[8][315] = 1;
   assign ecchmatrix[9][315] = 1;
   assign ecchmatrix[0][316] = 0;
   assign ecchmatrix[1][316] = 0;
   assign ecchmatrix[2][316] = 1;
   assign ecchmatrix[3][316] = 1;
   assign ecchmatrix[4][316] = 1;
   assign ecchmatrix[5][316] = 1;
   assign ecchmatrix[6][316] = 1;
   assign ecchmatrix[7][316] = 0;
   assign ecchmatrix[8][316] = 0;
   assign ecchmatrix[9][316] = 0;
   assign ecchmatrix[0][317] = 0;
   assign ecchmatrix[1][317] = 0;
   assign ecchmatrix[2][317] = 1;
   assign ecchmatrix[3][317] = 1;
   assign ecchmatrix[4][317] = 1;
   assign ecchmatrix[5][317] = 1;
   assign ecchmatrix[6][317] = 0;
   assign ecchmatrix[7][317] = 1;
   assign ecchmatrix[8][317] = 0;
   assign ecchmatrix[9][317] = 0;
   assign ecchmatrix[0][318] = 0;
   assign ecchmatrix[1][318] = 0;
   assign ecchmatrix[2][318] = 1;
   assign ecchmatrix[3][318] = 1;
   assign ecchmatrix[4][318] = 1;
   assign ecchmatrix[5][318] = 1;
   assign ecchmatrix[6][318] = 0;
   assign ecchmatrix[7][318] = 0;
   assign ecchmatrix[8][318] = 1;
   assign ecchmatrix[9][318] = 0;
   assign ecchmatrix[0][319] = 0;
   assign ecchmatrix[1][319] = 0;
   assign ecchmatrix[2][319] = 1;
   assign ecchmatrix[3][319] = 1;
   assign ecchmatrix[4][319] = 1;
   assign ecchmatrix[5][319] = 1;
   assign ecchmatrix[6][319] = 0;
   assign ecchmatrix[7][319] = 0;
   assign ecchmatrix[8][319] = 0;
   assign ecchmatrix[9][319] = 1;
   assign ecchmatrix[0][320] = 0;
   assign ecchmatrix[1][320] = 0;
   assign ecchmatrix[2][320] = 1;
   assign ecchmatrix[3][320] = 1;
   assign ecchmatrix[4][320] = 1;
   assign ecchmatrix[5][320] = 0;
   assign ecchmatrix[6][320] = 1;
   assign ecchmatrix[7][320] = 1;
   assign ecchmatrix[8][320] = 0;
   assign ecchmatrix[9][320] = 0;
   assign ecchmatrix[0][321] = 0;
   assign ecchmatrix[1][321] = 0;
   assign ecchmatrix[2][321] = 1;
   assign ecchmatrix[3][321] = 1;
   assign ecchmatrix[4][321] = 1;
   assign ecchmatrix[5][321] = 0;
   assign ecchmatrix[6][321] = 1;
   assign ecchmatrix[7][321] = 0;
   assign ecchmatrix[8][321] = 1;
   assign ecchmatrix[9][321] = 0;
   assign ecchmatrix[0][322] = 0;
   assign ecchmatrix[1][322] = 0;
   assign ecchmatrix[2][322] = 1;
   assign ecchmatrix[3][322] = 1;
   assign ecchmatrix[4][322] = 1;
   assign ecchmatrix[5][322] = 0;
   assign ecchmatrix[6][322] = 1;
   assign ecchmatrix[7][322] = 0;
   assign ecchmatrix[8][322] = 0;
   assign ecchmatrix[9][322] = 1;
   assign ecchmatrix[0][323] = 0;
   assign ecchmatrix[1][323] = 0;
   assign ecchmatrix[2][323] = 1;
   assign ecchmatrix[3][323] = 1;
   assign ecchmatrix[4][323] = 1;
   assign ecchmatrix[5][323] = 0;
   assign ecchmatrix[6][323] = 0;
   assign ecchmatrix[7][323] = 1;
   assign ecchmatrix[8][323] = 1;
   assign ecchmatrix[9][323] = 0;
   assign ecchmatrix[0][324] = 0;
   assign ecchmatrix[1][324] = 0;
   assign ecchmatrix[2][324] = 1;
   assign ecchmatrix[3][324] = 1;
   assign ecchmatrix[4][324] = 1;
   assign ecchmatrix[5][324] = 0;
   assign ecchmatrix[6][324] = 0;
   assign ecchmatrix[7][324] = 1;
   assign ecchmatrix[8][324] = 0;
   assign ecchmatrix[9][324] = 1;
   assign ecchmatrix[0][325] = 0;
   assign ecchmatrix[1][325] = 0;
   assign ecchmatrix[2][325] = 1;
   assign ecchmatrix[3][325] = 1;
   assign ecchmatrix[4][325] = 1;
   assign ecchmatrix[5][325] = 0;
   assign ecchmatrix[6][325] = 0;
   assign ecchmatrix[7][325] = 0;
   assign ecchmatrix[8][325] = 1;
   assign ecchmatrix[9][325] = 1;
   assign ecchmatrix[0][326] = 0;
   assign ecchmatrix[1][326] = 0;
   assign ecchmatrix[2][326] = 1;
   assign ecchmatrix[3][326] = 1;
   assign ecchmatrix[4][326] = 0;
   assign ecchmatrix[5][326] = 1;
   assign ecchmatrix[6][326] = 1;
   assign ecchmatrix[7][326] = 1;
   assign ecchmatrix[8][326] = 0;
   assign ecchmatrix[9][326] = 0;
   assign ecchmatrix[0][327] = 0;
   assign ecchmatrix[1][327] = 0;
   assign ecchmatrix[2][327] = 1;
   assign ecchmatrix[3][327] = 1;
   assign ecchmatrix[4][327] = 0;
   assign ecchmatrix[5][327] = 1;
   assign ecchmatrix[6][327] = 1;
   assign ecchmatrix[7][327] = 0;
   assign ecchmatrix[8][327] = 1;
   assign ecchmatrix[9][327] = 0;
   assign ecchmatrix[0][328] = 0;
   assign ecchmatrix[1][328] = 0;
   assign ecchmatrix[2][328] = 1;
   assign ecchmatrix[3][328] = 1;
   assign ecchmatrix[4][328] = 0;
   assign ecchmatrix[5][328] = 1;
   assign ecchmatrix[6][328] = 1;
   assign ecchmatrix[7][328] = 0;
   assign ecchmatrix[8][328] = 0;
   assign ecchmatrix[9][328] = 1;
   assign ecchmatrix[0][329] = 0;
   assign ecchmatrix[1][329] = 0;
   assign ecchmatrix[2][329] = 1;
   assign ecchmatrix[3][329] = 1;
   assign ecchmatrix[4][329] = 0;
   assign ecchmatrix[5][329] = 1;
   assign ecchmatrix[6][329] = 0;
   assign ecchmatrix[7][329] = 1;
   assign ecchmatrix[8][329] = 1;
   assign ecchmatrix[9][329] = 0;
   assign ecchmatrix[0][330] = 0;
   assign ecchmatrix[1][330] = 0;
   assign ecchmatrix[2][330] = 1;
   assign ecchmatrix[3][330] = 1;
   assign ecchmatrix[4][330] = 0;
   assign ecchmatrix[5][330] = 1;
   assign ecchmatrix[6][330] = 0;
   assign ecchmatrix[7][330] = 1;
   assign ecchmatrix[8][330] = 0;
   assign ecchmatrix[9][330] = 1;
   assign ecchmatrix[0][331] = 0;
   assign ecchmatrix[1][331] = 0;
   assign ecchmatrix[2][331] = 1;
   assign ecchmatrix[3][331] = 1;
   assign ecchmatrix[4][331] = 0;
   assign ecchmatrix[5][331] = 1;
   assign ecchmatrix[6][331] = 0;
   assign ecchmatrix[7][331] = 0;
   assign ecchmatrix[8][331] = 1;
   assign ecchmatrix[9][331] = 1;
   assign ecchmatrix[0][332] = 0;
   assign ecchmatrix[1][332] = 0;
   assign ecchmatrix[2][332] = 1;
   assign ecchmatrix[3][332] = 1;
   assign ecchmatrix[4][332] = 0;
   assign ecchmatrix[5][332] = 0;
   assign ecchmatrix[6][332] = 1;
   assign ecchmatrix[7][332] = 1;
   assign ecchmatrix[8][332] = 1;
   assign ecchmatrix[9][332] = 0;
   assign ecchmatrix[0][333] = 0;
   assign ecchmatrix[1][333] = 0;
   assign ecchmatrix[2][333] = 1;
   assign ecchmatrix[3][333] = 1;
   assign ecchmatrix[4][333] = 0;
   assign ecchmatrix[5][333] = 0;
   assign ecchmatrix[6][333] = 1;
   assign ecchmatrix[7][333] = 1;
   assign ecchmatrix[8][333] = 0;
   assign ecchmatrix[9][333] = 1;
   assign ecchmatrix[0][334] = 0;
   assign ecchmatrix[1][334] = 0;
   assign ecchmatrix[2][334] = 1;
   assign ecchmatrix[3][334] = 1;
   assign ecchmatrix[4][334] = 0;
   assign ecchmatrix[5][334] = 0;
   assign ecchmatrix[6][334] = 1;
   assign ecchmatrix[7][334] = 0;
   assign ecchmatrix[8][334] = 1;
   assign ecchmatrix[9][334] = 1;
   assign ecchmatrix[0][335] = 0;
   assign ecchmatrix[1][335] = 0;
   assign ecchmatrix[2][335] = 1;
   assign ecchmatrix[3][335] = 1;
   assign ecchmatrix[4][335] = 0;
   assign ecchmatrix[5][335] = 0;
   assign ecchmatrix[6][335] = 0;
   assign ecchmatrix[7][335] = 1;
   assign ecchmatrix[8][335] = 1;
   assign ecchmatrix[9][335] = 1;
   assign ecchmatrix[0][336] = 0;
   assign ecchmatrix[1][336] = 0;
   assign ecchmatrix[2][336] = 1;
   assign ecchmatrix[3][336] = 0;
   assign ecchmatrix[4][336] = 1;
   assign ecchmatrix[5][336] = 1;
   assign ecchmatrix[6][336] = 1;
   assign ecchmatrix[7][336] = 1;
   assign ecchmatrix[8][336] = 0;
   assign ecchmatrix[9][336] = 0;
   assign ecchmatrix[0][337] = 0;
   assign ecchmatrix[1][337] = 0;
   assign ecchmatrix[2][337] = 1;
   assign ecchmatrix[3][337] = 0;
   assign ecchmatrix[4][337] = 1;
   assign ecchmatrix[5][337] = 1;
   assign ecchmatrix[6][337] = 1;
   assign ecchmatrix[7][337] = 0;
   assign ecchmatrix[8][337] = 1;
   assign ecchmatrix[9][337] = 0;
   assign ecchmatrix[0][338] = 0;
   assign ecchmatrix[1][338] = 0;
   assign ecchmatrix[2][338] = 1;
   assign ecchmatrix[3][338] = 0;
   assign ecchmatrix[4][338] = 1;
   assign ecchmatrix[5][338] = 1;
   assign ecchmatrix[6][338] = 1;
   assign ecchmatrix[7][338] = 0;
   assign ecchmatrix[8][338] = 0;
   assign ecchmatrix[9][338] = 1;
   assign ecchmatrix[0][339] = 0;
   assign ecchmatrix[1][339] = 0;
   assign ecchmatrix[2][339] = 1;
   assign ecchmatrix[3][339] = 0;
   assign ecchmatrix[4][339] = 1;
   assign ecchmatrix[5][339] = 1;
   assign ecchmatrix[6][339] = 0;
   assign ecchmatrix[7][339] = 1;
   assign ecchmatrix[8][339] = 1;
   assign ecchmatrix[9][339] = 0;
   assign ecchmatrix[0][340] = 0;
   assign ecchmatrix[1][340] = 0;
   assign ecchmatrix[2][340] = 1;
   assign ecchmatrix[3][340] = 0;
   assign ecchmatrix[4][340] = 1;
   assign ecchmatrix[5][340] = 1;
   assign ecchmatrix[6][340] = 0;
   assign ecchmatrix[7][340] = 1;
   assign ecchmatrix[8][340] = 0;
   assign ecchmatrix[9][340] = 1;
   assign ecchmatrix[0][341] = 0;
   assign ecchmatrix[1][341] = 0;
   assign ecchmatrix[2][341] = 1;
   assign ecchmatrix[3][341] = 0;
   assign ecchmatrix[4][341] = 1;
   assign ecchmatrix[5][341] = 1;
   assign ecchmatrix[6][341] = 0;
   assign ecchmatrix[7][341] = 0;
   assign ecchmatrix[8][341] = 1;
   assign ecchmatrix[9][341] = 1;
   assign ecchmatrix[0][342] = 0;
   assign ecchmatrix[1][342] = 0;
   assign ecchmatrix[2][342] = 1;
   assign ecchmatrix[3][342] = 0;
   assign ecchmatrix[4][342] = 1;
   assign ecchmatrix[5][342] = 0;
   assign ecchmatrix[6][342] = 1;
   assign ecchmatrix[7][342] = 1;
   assign ecchmatrix[8][342] = 1;
   assign ecchmatrix[9][342] = 0;
   assign ecchmatrix[0][343] = 0;
   assign ecchmatrix[1][343] = 0;
   assign ecchmatrix[2][343] = 1;
   assign ecchmatrix[3][343] = 0;
   assign ecchmatrix[4][343] = 1;
   assign ecchmatrix[5][343] = 0;
   assign ecchmatrix[6][343] = 1;
   assign ecchmatrix[7][343] = 1;
   assign ecchmatrix[8][343] = 0;
   assign ecchmatrix[9][343] = 1;
   assign ecchmatrix[0][344] = 0;
   assign ecchmatrix[1][344] = 0;
   assign ecchmatrix[2][344] = 1;
   assign ecchmatrix[3][344] = 0;
   assign ecchmatrix[4][344] = 1;
   assign ecchmatrix[5][344] = 0;
   assign ecchmatrix[6][344] = 1;
   assign ecchmatrix[7][344] = 0;
   assign ecchmatrix[8][344] = 1;
   assign ecchmatrix[9][344] = 1;
   assign ecchmatrix[0][345] = 0;
   assign ecchmatrix[1][345] = 0;
   assign ecchmatrix[2][345] = 1;
   assign ecchmatrix[3][345] = 0;
   assign ecchmatrix[4][345] = 1;
   assign ecchmatrix[5][345] = 0;
   assign ecchmatrix[6][345] = 0;
   assign ecchmatrix[7][345] = 1;
   assign ecchmatrix[8][345] = 1;
   assign ecchmatrix[9][345] = 1;
   assign ecchmatrix[0][346] = 0;
   assign ecchmatrix[1][346] = 0;
   assign ecchmatrix[2][346] = 1;
   assign ecchmatrix[3][346] = 0;
   assign ecchmatrix[4][346] = 0;
   assign ecchmatrix[5][346] = 1;
   assign ecchmatrix[6][346] = 1;
   assign ecchmatrix[7][346] = 1;
   assign ecchmatrix[8][346] = 1;
   assign ecchmatrix[9][346] = 0;
   assign ecchmatrix[0][347] = 0;
   assign ecchmatrix[1][347] = 0;
   assign ecchmatrix[2][347] = 1;
   assign ecchmatrix[3][347] = 0;
   assign ecchmatrix[4][347] = 0;
   assign ecchmatrix[5][347] = 1;
   assign ecchmatrix[6][347] = 1;
   assign ecchmatrix[7][347] = 1;
   assign ecchmatrix[8][347] = 0;
   assign ecchmatrix[9][347] = 1;
   assign ecchmatrix[0][348] = 0;
   assign ecchmatrix[1][348] = 0;
   assign ecchmatrix[2][348] = 1;
   assign ecchmatrix[3][348] = 0;
   assign ecchmatrix[4][348] = 0;
   assign ecchmatrix[5][348] = 1;
   assign ecchmatrix[6][348] = 1;
   assign ecchmatrix[7][348] = 0;
   assign ecchmatrix[8][348] = 1;
   assign ecchmatrix[9][348] = 1;
   assign ecchmatrix[0][349] = 0;
   assign ecchmatrix[1][349] = 0;
   assign ecchmatrix[2][349] = 1;
   assign ecchmatrix[3][349] = 0;
   assign ecchmatrix[4][349] = 0;
   assign ecchmatrix[5][349] = 1;
   assign ecchmatrix[6][349] = 0;
   assign ecchmatrix[7][349] = 1;
   assign ecchmatrix[8][349] = 1;
   assign ecchmatrix[9][349] = 1;
   assign ecchmatrix[0][350] = 0;
   assign ecchmatrix[1][350] = 0;
   assign ecchmatrix[2][350] = 1;
   assign ecchmatrix[3][350] = 0;
   assign ecchmatrix[4][350] = 0;
   assign ecchmatrix[5][350] = 0;
   assign ecchmatrix[6][350] = 1;
   assign ecchmatrix[7][350] = 1;
   assign ecchmatrix[8][350] = 1;
   assign ecchmatrix[9][350] = 1;
   assign ecchmatrix[0][351] = 0;
   assign ecchmatrix[1][351] = 0;
   assign ecchmatrix[2][351] = 0;
   assign ecchmatrix[3][351] = 1;
   assign ecchmatrix[4][351] = 1;
   assign ecchmatrix[5][351] = 1;
   assign ecchmatrix[6][351] = 1;
   assign ecchmatrix[7][351] = 1;
   assign ecchmatrix[8][351] = 0;
   assign ecchmatrix[9][351] = 0;
   assign ecchmatrix[0][352] = 0;
   assign ecchmatrix[1][352] = 0;
   assign ecchmatrix[2][352] = 0;
   assign ecchmatrix[3][352] = 1;
   assign ecchmatrix[4][352] = 1;
   assign ecchmatrix[5][352] = 1;
   assign ecchmatrix[6][352] = 1;
   assign ecchmatrix[7][352] = 0;
   assign ecchmatrix[8][352] = 1;
   assign ecchmatrix[9][352] = 0;
   assign ecchmatrix[0][353] = 0;
   assign ecchmatrix[1][353] = 0;
   assign ecchmatrix[2][353] = 0;
   assign ecchmatrix[3][353] = 1;
   assign ecchmatrix[4][353] = 1;
   assign ecchmatrix[5][353] = 1;
   assign ecchmatrix[6][353] = 1;
   assign ecchmatrix[7][353] = 0;
   assign ecchmatrix[8][353] = 0;
   assign ecchmatrix[9][353] = 1;
   assign ecchmatrix[0][354] = 0;
   assign ecchmatrix[1][354] = 0;
   assign ecchmatrix[2][354] = 0;
   assign ecchmatrix[3][354] = 1;
   assign ecchmatrix[4][354] = 1;
   assign ecchmatrix[5][354] = 1;
   assign ecchmatrix[6][354] = 0;
   assign ecchmatrix[7][354] = 1;
   assign ecchmatrix[8][354] = 1;
   assign ecchmatrix[9][354] = 0;
   assign ecchmatrix[0][355] = 0;
   assign ecchmatrix[1][355] = 0;
   assign ecchmatrix[2][355] = 0;
   assign ecchmatrix[3][355] = 1;
   assign ecchmatrix[4][355] = 1;
   assign ecchmatrix[5][355] = 1;
   assign ecchmatrix[6][355] = 0;
   assign ecchmatrix[7][355] = 1;
   assign ecchmatrix[8][355] = 0;
   assign ecchmatrix[9][355] = 1;
   assign ecchmatrix[0][356] = 0;
   assign ecchmatrix[1][356] = 0;
   assign ecchmatrix[2][356] = 0;
   assign ecchmatrix[3][356] = 1;
   assign ecchmatrix[4][356] = 1;
   assign ecchmatrix[5][356] = 1;
   assign ecchmatrix[6][356] = 0;
   assign ecchmatrix[7][356] = 0;
   assign ecchmatrix[8][356] = 1;
   assign ecchmatrix[9][356] = 1;
   assign ecchmatrix[0][357] = 0;
   assign ecchmatrix[1][357] = 0;
   assign ecchmatrix[2][357] = 0;
   assign ecchmatrix[3][357] = 1;
   assign ecchmatrix[4][357] = 1;
   assign ecchmatrix[5][357] = 0;
   assign ecchmatrix[6][357] = 1;
   assign ecchmatrix[7][357] = 1;
   assign ecchmatrix[8][357] = 1;
   assign ecchmatrix[9][357] = 0;
   assign ecchmatrix[0][358] = 0;
   assign ecchmatrix[1][358] = 0;
   assign ecchmatrix[2][358] = 0;
   assign ecchmatrix[3][358] = 1;
   assign ecchmatrix[4][358] = 1;
   assign ecchmatrix[5][358] = 0;
   assign ecchmatrix[6][358] = 1;
   assign ecchmatrix[7][358] = 1;
   assign ecchmatrix[8][358] = 0;
   assign ecchmatrix[9][358] = 1;
   assign ecchmatrix[0][359] = 0;
   assign ecchmatrix[1][359] = 0;
   assign ecchmatrix[2][359] = 0;
   assign ecchmatrix[3][359] = 1;
   assign ecchmatrix[4][359] = 1;
   assign ecchmatrix[5][359] = 0;
   assign ecchmatrix[6][359] = 1;
   assign ecchmatrix[7][359] = 0;
   assign ecchmatrix[8][359] = 1;
   assign ecchmatrix[9][359] = 1;
   assign ecchmatrix[0][360] = 0;
   assign ecchmatrix[1][360] = 0;
   assign ecchmatrix[2][360] = 0;
   assign ecchmatrix[3][360] = 1;
   assign ecchmatrix[4][360] = 1;
   assign ecchmatrix[5][360] = 0;
   assign ecchmatrix[6][360] = 0;
   assign ecchmatrix[7][360] = 1;
   assign ecchmatrix[8][360] = 1;
   assign ecchmatrix[9][360] = 1;
   assign ecchmatrix[0][361] = 0;
   assign ecchmatrix[1][361] = 0;
   assign ecchmatrix[2][361] = 0;
   assign ecchmatrix[3][361] = 1;
   assign ecchmatrix[4][361] = 0;
   assign ecchmatrix[5][361] = 1;
   assign ecchmatrix[6][361] = 1;
   assign ecchmatrix[7][361] = 1;
   assign ecchmatrix[8][361] = 1;
   assign ecchmatrix[9][361] = 0;
   assign ecchmatrix[0][362] = 0;
   assign ecchmatrix[1][362] = 0;
   assign ecchmatrix[2][362] = 0;
   assign ecchmatrix[3][362] = 1;
   assign ecchmatrix[4][362] = 0;
   assign ecchmatrix[5][362] = 1;
   assign ecchmatrix[6][362] = 1;
   assign ecchmatrix[7][362] = 1;
   assign ecchmatrix[8][362] = 0;
   assign ecchmatrix[9][362] = 1;
   assign ecchmatrix[0][363] = 0;
   assign ecchmatrix[1][363] = 0;
   assign ecchmatrix[2][363] = 0;
   assign ecchmatrix[3][363] = 1;
   assign ecchmatrix[4][363] = 0;
   assign ecchmatrix[5][363] = 1;
   assign ecchmatrix[6][363] = 1;
   assign ecchmatrix[7][363] = 0;
   assign ecchmatrix[8][363] = 1;
   assign ecchmatrix[9][363] = 1;
   assign ecchmatrix[0][364] = 0;
   assign ecchmatrix[1][364] = 0;
   assign ecchmatrix[2][364] = 0;
   assign ecchmatrix[3][364] = 1;
   assign ecchmatrix[4][364] = 0;
   assign ecchmatrix[5][364] = 1;
   assign ecchmatrix[6][364] = 0;
   assign ecchmatrix[7][364] = 1;
   assign ecchmatrix[8][364] = 1;
   assign ecchmatrix[9][364] = 1;
   assign ecchmatrix[0][365] = 0;
   assign ecchmatrix[1][365] = 0;
   assign ecchmatrix[2][365] = 0;
   assign ecchmatrix[3][365] = 1;
   assign ecchmatrix[4][365] = 0;
   assign ecchmatrix[5][365] = 0;
   assign ecchmatrix[6][365] = 1;
   assign ecchmatrix[7][365] = 1;
   assign ecchmatrix[8][365] = 1;
   assign ecchmatrix[9][365] = 1;
   assign ecchmatrix[0][366] = 0;
   assign ecchmatrix[1][366] = 0;
   assign ecchmatrix[2][366] = 0;
   assign ecchmatrix[3][366] = 0;
   assign ecchmatrix[4][366] = 1;
   assign ecchmatrix[5][366] = 1;
   assign ecchmatrix[6][366] = 1;
   assign ecchmatrix[7][366] = 1;
   assign ecchmatrix[8][366] = 1;
   assign ecchmatrix[9][366] = 0;
   assign ecchmatrix[0][367] = 0;
   assign ecchmatrix[1][367] = 0;
   assign ecchmatrix[2][367] = 0;
   assign ecchmatrix[3][367] = 0;
   assign ecchmatrix[4][367] = 1;
   assign ecchmatrix[5][367] = 1;
   assign ecchmatrix[6][367] = 1;
   assign ecchmatrix[7][367] = 1;
   assign ecchmatrix[8][367] = 0;
   assign ecchmatrix[9][367] = 1;
   assign ecchmatrix[0][368] = 0;
   assign ecchmatrix[1][368] = 0;
   assign ecchmatrix[2][368] = 0;
   assign ecchmatrix[3][368] = 0;
   assign ecchmatrix[4][368] = 1;
   assign ecchmatrix[5][368] = 1;
   assign ecchmatrix[6][368] = 1;
   assign ecchmatrix[7][368] = 0;
   assign ecchmatrix[8][368] = 1;
   assign ecchmatrix[9][368] = 1;
   assign ecchmatrix[0][369] = 0;
   assign ecchmatrix[1][369] = 0;
   assign ecchmatrix[2][369] = 0;
   assign ecchmatrix[3][369] = 0;
   assign ecchmatrix[4][369] = 1;
   assign ecchmatrix[5][369] = 1;
   assign ecchmatrix[6][369] = 0;
   assign ecchmatrix[7][369] = 1;
   assign ecchmatrix[8][369] = 1;
   assign ecchmatrix[9][369] = 1;
   assign ecchmatrix[0][370] = 0;
   assign ecchmatrix[1][370] = 0;
   assign ecchmatrix[2][370] = 0;
   assign ecchmatrix[3][370] = 0;
   assign ecchmatrix[4][370] = 1;
   assign ecchmatrix[5][370] = 0;
   assign ecchmatrix[6][370] = 1;
   assign ecchmatrix[7][370] = 1;
   assign ecchmatrix[8][370] = 1;
   assign ecchmatrix[9][370] = 1;
   assign ecchmatrix[0][371] = 0;
   assign ecchmatrix[1][371] = 0;
   assign ecchmatrix[2][371] = 0;
   assign ecchmatrix[3][371] = 0;
   assign ecchmatrix[4][371] = 0;
   assign ecchmatrix[5][371] = 1;
   assign ecchmatrix[6][371] = 1;
   assign ecchmatrix[7][371] = 1;
   assign ecchmatrix[8][371] = 1;
   assign ecchmatrix[9][371] = 1;
   assign ecchmatrix[0][372] = 1;
   assign ecchmatrix[1][372] = 1;
   assign ecchmatrix[2][372] = 1;
   assign ecchmatrix[3][372] = 1;
   assign ecchmatrix[4][372] = 1;
   assign ecchmatrix[5][372] = 1;
   assign ecchmatrix[6][372] = 1;
   assign ecchmatrix[7][372] = 0;
   assign ecchmatrix[8][372] = 0;
   assign ecchmatrix[9][372] = 0;
   assign ecchmatrix[0][373] = 1;
   assign ecchmatrix[1][373] = 1;
   assign ecchmatrix[2][373] = 1;
   assign ecchmatrix[3][373] = 1;
   assign ecchmatrix[4][373] = 1;
   assign ecchmatrix[5][373] = 1;
   assign ecchmatrix[6][373] = 0;
   assign ecchmatrix[7][373] = 1;
   assign ecchmatrix[8][373] = 0;
   assign ecchmatrix[9][373] = 0;
   assign ecchmatrix[0][374] = 1;
   assign ecchmatrix[1][374] = 1;
   assign ecchmatrix[2][374] = 1;
   assign ecchmatrix[3][374] = 1;
   assign ecchmatrix[4][374] = 1;
   assign ecchmatrix[5][374] = 1;
   assign ecchmatrix[6][374] = 0;
   assign ecchmatrix[7][374] = 0;
   assign ecchmatrix[8][374] = 1;
   assign ecchmatrix[9][374] = 0;
   assign ecchmatrix[0][375] = 1;
   assign ecchmatrix[1][375] = 1;
   assign ecchmatrix[2][375] = 1;
   assign ecchmatrix[3][375] = 1;
   assign ecchmatrix[4][375] = 1;
   assign ecchmatrix[5][375] = 1;
   assign ecchmatrix[6][375] = 0;
   assign ecchmatrix[7][375] = 0;
   assign ecchmatrix[8][375] = 0;
   assign ecchmatrix[9][375] = 1;
   assign ecchmatrix[0][376] = 1;
   assign ecchmatrix[1][376] = 1;
   assign ecchmatrix[2][376] = 1;
   assign ecchmatrix[3][376] = 1;
   assign ecchmatrix[4][376] = 1;
   assign ecchmatrix[5][376] = 0;
   assign ecchmatrix[6][376] = 1;
   assign ecchmatrix[7][376] = 1;
   assign ecchmatrix[8][376] = 0;
   assign ecchmatrix[9][376] = 0;
   assign ecchmatrix[0][377] = 1;
   assign ecchmatrix[1][377] = 1;
   assign ecchmatrix[2][377] = 1;
   assign ecchmatrix[3][377] = 1;
   assign ecchmatrix[4][377] = 1;
   assign ecchmatrix[5][377] = 0;
   assign ecchmatrix[6][377] = 1;
   assign ecchmatrix[7][377] = 0;
   assign ecchmatrix[8][377] = 1;
   assign ecchmatrix[9][377] = 0;
   assign ecchmatrix[0][378] = 1;
   assign ecchmatrix[1][378] = 1;
   assign ecchmatrix[2][378] = 1;
   assign ecchmatrix[3][378] = 1;
   assign ecchmatrix[4][378] = 1;
   assign ecchmatrix[5][378] = 0;
   assign ecchmatrix[6][378] = 1;
   assign ecchmatrix[7][378] = 0;
   assign ecchmatrix[8][378] = 0;
   assign ecchmatrix[9][378] = 1;
   assign ecchmatrix[0][379] = 1;
   assign ecchmatrix[1][379] = 1;
   assign ecchmatrix[2][379] = 1;
   assign ecchmatrix[3][379] = 1;
   assign ecchmatrix[4][379] = 1;
   assign ecchmatrix[5][379] = 0;
   assign ecchmatrix[6][379] = 0;
   assign ecchmatrix[7][379] = 1;
   assign ecchmatrix[8][379] = 1;
   assign ecchmatrix[9][379] = 0;
   assign ecchmatrix[0][380] = 1;
   assign ecchmatrix[1][380] = 1;
   assign ecchmatrix[2][380] = 1;
   assign ecchmatrix[3][380] = 1;
   assign ecchmatrix[4][380] = 1;
   assign ecchmatrix[5][380] = 0;
   assign ecchmatrix[6][380] = 0;
   assign ecchmatrix[7][380] = 1;
   assign ecchmatrix[8][380] = 0;
   assign ecchmatrix[9][380] = 1;
   assign ecchmatrix[0][381] = 1;
   assign ecchmatrix[1][381] = 1;
   assign ecchmatrix[2][381] = 1;
   assign ecchmatrix[3][381] = 1;
   assign ecchmatrix[4][381] = 1;
   assign ecchmatrix[5][381] = 0;
   assign ecchmatrix[6][381] = 0;
   assign ecchmatrix[7][381] = 0;
   assign ecchmatrix[8][381] = 1;
   assign ecchmatrix[9][381] = 1;
   assign ecchmatrix[0][382] = 1;
   assign ecchmatrix[1][382] = 1;
   assign ecchmatrix[2][382] = 1;
   assign ecchmatrix[3][382] = 1;
   assign ecchmatrix[4][382] = 0;
   assign ecchmatrix[5][382] = 1;
   assign ecchmatrix[6][382] = 1;
   assign ecchmatrix[7][382] = 1;
   assign ecchmatrix[8][382] = 0;
   assign ecchmatrix[9][382] = 0;
   assign ecchmatrix[0][383] = 1;
   assign ecchmatrix[1][383] = 1;
   assign ecchmatrix[2][383] = 1;
   assign ecchmatrix[3][383] = 1;
   assign ecchmatrix[4][383] = 0;
   assign ecchmatrix[5][383] = 1;
   assign ecchmatrix[6][383] = 1;
   assign ecchmatrix[7][383] = 0;
   assign ecchmatrix[8][383] = 1;
   assign ecchmatrix[9][383] = 0;
   assign ecchmatrix[0][384] = 1;
   assign ecchmatrix[1][384] = 1;
   assign ecchmatrix[2][384] = 1;
   assign ecchmatrix[3][384] = 1;
   assign ecchmatrix[4][384] = 0;
   assign ecchmatrix[5][384] = 1;
   assign ecchmatrix[6][384] = 1;
   assign ecchmatrix[7][384] = 0;
   assign ecchmatrix[8][384] = 0;
   assign ecchmatrix[9][384] = 1;
   assign ecchmatrix[0][385] = 1;
   assign ecchmatrix[1][385] = 1;
   assign ecchmatrix[2][385] = 1;
   assign ecchmatrix[3][385] = 1;
   assign ecchmatrix[4][385] = 0;
   assign ecchmatrix[5][385] = 1;
   assign ecchmatrix[6][385] = 0;
   assign ecchmatrix[7][385] = 1;
   assign ecchmatrix[8][385] = 1;
   assign ecchmatrix[9][385] = 0;
   assign ecchmatrix[0][386] = 1;
   assign ecchmatrix[1][386] = 1;
   assign ecchmatrix[2][386] = 1;
   assign ecchmatrix[3][386] = 1;
   assign ecchmatrix[4][386] = 0;
   assign ecchmatrix[5][386] = 1;
   assign ecchmatrix[6][386] = 0;
   assign ecchmatrix[7][386] = 1;
   assign ecchmatrix[8][386] = 0;
   assign ecchmatrix[9][386] = 1;
   assign ecchmatrix[0][387] = 1;
   assign ecchmatrix[1][387] = 1;
   assign ecchmatrix[2][387] = 1;
   assign ecchmatrix[3][387] = 1;
   assign ecchmatrix[4][387] = 0;
   assign ecchmatrix[5][387] = 1;
   assign ecchmatrix[6][387] = 0;
   assign ecchmatrix[7][387] = 0;
   assign ecchmatrix[8][387] = 1;
   assign ecchmatrix[9][387] = 1;
   assign ecchmatrix[0][388] = 1;
   assign ecchmatrix[1][388] = 1;
   assign ecchmatrix[2][388] = 1;
   assign ecchmatrix[3][388] = 1;
   assign ecchmatrix[4][388] = 0;
   assign ecchmatrix[5][388] = 0;
   assign ecchmatrix[6][388] = 1;
   assign ecchmatrix[7][388] = 1;
   assign ecchmatrix[8][388] = 1;
   assign ecchmatrix[9][388] = 0;
   assign ecchmatrix[0][389] = 1;
   assign ecchmatrix[1][389] = 1;
   assign ecchmatrix[2][389] = 1;
   assign ecchmatrix[3][389] = 1;
   assign ecchmatrix[4][389] = 0;
   assign ecchmatrix[5][389] = 0;
   assign ecchmatrix[6][389] = 1;
   assign ecchmatrix[7][389] = 1;
   assign ecchmatrix[8][389] = 0;
   assign ecchmatrix[9][389] = 1;
   assign ecchmatrix[0][390] = 1;
   assign ecchmatrix[1][390] = 1;
   assign ecchmatrix[2][390] = 1;
   assign ecchmatrix[3][390] = 1;
   assign ecchmatrix[4][390] = 0;
   assign ecchmatrix[5][390] = 0;
   assign ecchmatrix[6][390] = 1;
   assign ecchmatrix[7][390] = 0;
   assign ecchmatrix[8][390] = 1;
   assign ecchmatrix[9][390] = 1;
   assign ecchmatrix[0][391] = 1;
   assign ecchmatrix[1][391] = 1;
   assign ecchmatrix[2][391] = 1;
   assign ecchmatrix[3][391] = 1;
   assign ecchmatrix[4][391] = 0;
   assign ecchmatrix[5][391] = 0;
   assign ecchmatrix[6][391] = 0;
   assign ecchmatrix[7][391] = 1;
   assign ecchmatrix[8][391] = 1;
   assign ecchmatrix[9][391] = 1;
   assign ecchmatrix[0][392] = 1;
   assign ecchmatrix[1][392] = 1;
   assign ecchmatrix[2][392] = 1;
   assign ecchmatrix[3][392] = 0;
   assign ecchmatrix[4][392] = 1;
   assign ecchmatrix[5][392] = 1;
   assign ecchmatrix[6][392] = 1;
   assign ecchmatrix[7][392] = 1;
   assign ecchmatrix[8][392] = 0;
   assign ecchmatrix[9][392] = 0;
   assign ecchmatrix[0][393] = 1;
   assign ecchmatrix[1][393] = 1;
   assign ecchmatrix[2][393] = 1;
   assign ecchmatrix[3][393] = 0;
   assign ecchmatrix[4][393] = 1;
   assign ecchmatrix[5][393] = 1;
   assign ecchmatrix[6][393] = 1;
   assign ecchmatrix[7][393] = 0;
   assign ecchmatrix[8][393] = 1;
   assign ecchmatrix[9][393] = 0;
   assign ecchmatrix[0][394] = 1;
   assign ecchmatrix[1][394] = 1;
   assign ecchmatrix[2][394] = 1;
   assign ecchmatrix[3][394] = 0;
   assign ecchmatrix[4][394] = 1;
   assign ecchmatrix[5][394] = 1;
   assign ecchmatrix[6][394] = 1;
   assign ecchmatrix[7][394] = 0;
   assign ecchmatrix[8][394] = 0;
   assign ecchmatrix[9][394] = 1;
   assign ecchmatrix[0][395] = 1;
   assign ecchmatrix[1][395] = 1;
   assign ecchmatrix[2][395] = 1;
   assign ecchmatrix[3][395] = 0;
   assign ecchmatrix[4][395] = 1;
   assign ecchmatrix[5][395] = 1;
   assign ecchmatrix[6][395] = 0;
   assign ecchmatrix[7][395] = 1;
   assign ecchmatrix[8][395] = 1;
   assign ecchmatrix[9][395] = 0;
   assign ecchmatrix[0][396] = 1;
   assign ecchmatrix[1][396] = 1;
   assign ecchmatrix[2][396] = 1;
   assign ecchmatrix[3][396] = 0;
   assign ecchmatrix[4][396] = 1;
   assign ecchmatrix[5][396] = 1;
   assign ecchmatrix[6][396] = 0;
   assign ecchmatrix[7][396] = 1;
   assign ecchmatrix[8][396] = 0;
   assign ecchmatrix[9][396] = 1;
   assign ecchmatrix[0][397] = 1;
   assign ecchmatrix[1][397] = 1;
   assign ecchmatrix[2][397] = 1;
   assign ecchmatrix[3][397] = 0;
   assign ecchmatrix[4][397] = 1;
   assign ecchmatrix[5][397] = 1;
   assign ecchmatrix[6][397] = 0;
   assign ecchmatrix[7][397] = 0;
   assign ecchmatrix[8][397] = 1;
   assign ecchmatrix[9][397] = 1;
   assign ecchmatrix[0][398] = 1;
   assign ecchmatrix[1][398] = 1;
   assign ecchmatrix[2][398] = 1;
   assign ecchmatrix[3][398] = 0;
   assign ecchmatrix[4][398] = 1;
   assign ecchmatrix[5][398] = 0;
   assign ecchmatrix[6][398] = 1;
   assign ecchmatrix[7][398] = 1;
   assign ecchmatrix[8][398] = 1;
   assign ecchmatrix[9][398] = 0;
   assign ecchmatrix[0][399] = 1;
   assign ecchmatrix[1][399] = 1;
   assign ecchmatrix[2][399] = 1;
   assign ecchmatrix[3][399] = 0;
   assign ecchmatrix[4][399] = 1;
   assign ecchmatrix[5][399] = 0;
   assign ecchmatrix[6][399] = 1;
   assign ecchmatrix[7][399] = 1;
   assign ecchmatrix[8][399] = 0;
   assign ecchmatrix[9][399] = 1;
   assign ecchmatrix[0][400] = 1;
   assign ecchmatrix[1][400] = 1;
   assign ecchmatrix[2][400] = 1;
   assign ecchmatrix[3][400] = 0;
   assign ecchmatrix[4][400] = 1;
   assign ecchmatrix[5][400] = 0;
   assign ecchmatrix[6][400] = 1;
   assign ecchmatrix[7][400] = 0;
   assign ecchmatrix[8][400] = 1;
   assign ecchmatrix[9][400] = 1;
   assign ecchmatrix[0][401] = 1;
   assign ecchmatrix[1][401] = 1;
   assign ecchmatrix[2][401] = 1;
   assign ecchmatrix[3][401] = 0;
   assign ecchmatrix[4][401] = 1;
   assign ecchmatrix[5][401] = 0;
   assign ecchmatrix[6][401] = 0;
   assign ecchmatrix[7][401] = 1;
   assign ecchmatrix[8][401] = 1;
   assign ecchmatrix[9][401] = 1;
   assign ecchmatrix[0][402] = 1;
   assign ecchmatrix[1][402] = 1;
   assign ecchmatrix[2][402] = 1;
   assign ecchmatrix[3][402] = 0;
   assign ecchmatrix[4][402] = 0;
   assign ecchmatrix[5][402] = 1;
   assign ecchmatrix[6][402] = 1;
   assign ecchmatrix[7][402] = 1;
   assign ecchmatrix[8][402] = 1;
   assign ecchmatrix[9][402] = 0;
   assign ecchmatrix[0][403] = 1;
   assign ecchmatrix[1][403] = 1;
   assign ecchmatrix[2][403] = 1;
   assign ecchmatrix[3][403] = 0;
   assign ecchmatrix[4][403] = 0;
   assign ecchmatrix[5][403] = 1;
   assign ecchmatrix[6][403] = 1;
   assign ecchmatrix[7][403] = 1;
   assign ecchmatrix[8][403] = 0;
   assign ecchmatrix[9][403] = 1;
   assign ecchmatrix[0][404] = 1;
   assign ecchmatrix[1][404] = 1;
   assign ecchmatrix[2][404] = 1;
   assign ecchmatrix[3][404] = 0;
   assign ecchmatrix[4][404] = 0;
   assign ecchmatrix[5][404] = 1;
   assign ecchmatrix[6][404] = 1;
   assign ecchmatrix[7][404] = 0;
   assign ecchmatrix[8][404] = 1;
   assign ecchmatrix[9][404] = 1;
   assign ecchmatrix[0][405] = 1;
   assign ecchmatrix[1][405] = 1;
   assign ecchmatrix[2][405] = 1;
   assign ecchmatrix[3][405] = 0;
   assign ecchmatrix[4][405] = 0;
   assign ecchmatrix[5][405] = 1;
   assign ecchmatrix[6][405] = 0;
   assign ecchmatrix[7][405] = 1;
   assign ecchmatrix[8][405] = 1;
   assign ecchmatrix[9][405] = 1;
   assign ecchmatrix[0][406] = 1;
   assign ecchmatrix[1][406] = 1;
   assign ecchmatrix[2][406] = 1;
   assign ecchmatrix[3][406] = 0;
   assign ecchmatrix[4][406] = 0;
   assign ecchmatrix[5][406] = 0;
   assign ecchmatrix[6][406] = 1;
   assign ecchmatrix[7][406] = 1;
   assign ecchmatrix[8][406] = 1;
   assign ecchmatrix[9][406] = 1;
   assign ecchmatrix[0][407] = 1;
   assign ecchmatrix[1][407] = 1;
   assign ecchmatrix[2][407] = 0;
   assign ecchmatrix[3][407] = 1;
   assign ecchmatrix[4][407] = 1;
   assign ecchmatrix[5][407] = 1;
   assign ecchmatrix[6][407] = 1;
   assign ecchmatrix[7][407] = 1;
   assign ecchmatrix[8][407] = 0;
   assign ecchmatrix[9][407] = 0;
   assign ecchmatrix[0][408] = 1;
   assign ecchmatrix[1][408] = 1;
   assign ecchmatrix[2][408] = 0;
   assign ecchmatrix[3][408] = 1;
   assign ecchmatrix[4][408] = 1;
   assign ecchmatrix[5][408] = 1;
   assign ecchmatrix[6][408] = 1;
   assign ecchmatrix[7][408] = 0;
   assign ecchmatrix[8][408] = 1;
   assign ecchmatrix[9][408] = 0;
   assign ecchmatrix[0][409] = 1;
   assign ecchmatrix[1][409] = 1;
   assign ecchmatrix[2][409] = 0;
   assign ecchmatrix[3][409] = 1;
   assign ecchmatrix[4][409] = 1;
   assign ecchmatrix[5][409] = 1;
   assign ecchmatrix[6][409] = 1;
   assign ecchmatrix[7][409] = 0;
   assign ecchmatrix[8][409] = 0;
   assign ecchmatrix[9][409] = 1;
   assign ecchmatrix[0][410] = 1;
   assign ecchmatrix[1][410] = 1;
   assign ecchmatrix[2][410] = 0;
   assign ecchmatrix[3][410] = 1;
   assign ecchmatrix[4][410] = 1;
   assign ecchmatrix[5][410] = 1;
   assign ecchmatrix[6][410] = 0;
   assign ecchmatrix[7][410] = 1;
   assign ecchmatrix[8][410] = 1;
   assign ecchmatrix[9][410] = 0;
   assign ecchmatrix[0][411] = 1;
   assign ecchmatrix[1][411] = 1;
   assign ecchmatrix[2][411] = 0;
   assign ecchmatrix[3][411] = 1;
   assign ecchmatrix[4][411] = 1;
   assign ecchmatrix[5][411] = 1;
   assign ecchmatrix[6][411] = 0;
   assign ecchmatrix[7][411] = 1;
   assign ecchmatrix[8][411] = 0;
   assign ecchmatrix[9][411] = 1;
   assign ecchmatrix[0][412] = 1;
   assign ecchmatrix[1][412] = 1;
   assign ecchmatrix[2][412] = 0;
   assign ecchmatrix[3][412] = 1;
   assign ecchmatrix[4][412] = 1;
   assign ecchmatrix[5][412] = 1;
   assign ecchmatrix[6][412] = 0;
   assign ecchmatrix[7][412] = 0;
   assign ecchmatrix[8][412] = 1;
   assign ecchmatrix[9][412] = 1;
   assign ecchmatrix[0][413] = 1;
   assign ecchmatrix[1][413] = 1;
   assign ecchmatrix[2][413] = 0;
   assign ecchmatrix[3][413] = 1;
   assign ecchmatrix[4][413] = 1;
   assign ecchmatrix[5][413] = 0;
   assign ecchmatrix[6][413] = 1;
   assign ecchmatrix[7][413] = 1;
   assign ecchmatrix[8][413] = 1;
   assign ecchmatrix[9][413] = 0;
   assign ecchmatrix[0][414] = 1;
   assign ecchmatrix[1][414] = 1;
   assign ecchmatrix[2][414] = 0;
   assign ecchmatrix[3][414] = 1;
   assign ecchmatrix[4][414] = 1;
   assign ecchmatrix[5][414] = 0;
   assign ecchmatrix[6][414] = 1;
   assign ecchmatrix[7][414] = 1;
   assign ecchmatrix[8][414] = 0;
   assign ecchmatrix[9][414] = 1;
   assign ecchmatrix[0][415] = 1;
   assign ecchmatrix[1][415] = 1;
   assign ecchmatrix[2][415] = 0;
   assign ecchmatrix[3][415] = 1;
   assign ecchmatrix[4][415] = 1;
   assign ecchmatrix[5][415] = 0;
   assign ecchmatrix[6][415] = 1;
   assign ecchmatrix[7][415] = 0;
   assign ecchmatrix[8][415] = 1;
   assign ecchmatrix[9][415] = 1;
   assign ecchmatrix[0][416] = 1;
   assign ecchmatrix[1][416] = 1;
   assign ecchmatrix[2][416] = 0;
   assign ecchmatrix[3][416] = 1;
   assign ecchmatrix[4][416] = 1;
   assign ecchmatrix[5][416] = 0;
   assign ecchmatrix[6][416] = 0;
   assign ecchmatrix[7][416] = 1;
   assign ecchmatrix[8][416] = 1;
   assign ecchmatrix[9][416] = 1;
   assign ecchmatrix[0][417] = 1;
   assign ecchmatrix[1][417] = 1;
   assign ecchmatrix[2][417] = 0;
   assign ecchmatrix[3][417] = 1;
   assign ecchmatrix[4][417] = 0;
   assign ecchmatrix[5][417] = 1;
   assign ecchmatrix[6][417] = 1;
   assign ecchmatrix[7][417] = 1;
   assign ecchmatrix[8][417] = 1;
   assign ecchmatrix[9][417] = 0;
   assign ecchmatrix[0][418] = 1;
   assign ecchmatrix[1][418] = 1;
   assign ecchmatrix[2][418] = 0;
   assign ecchmatrix[3][418] = 1;
   assign ecchmatrix[4][418] = 0;
   assign ecchmatrix[5][418] = 1;
   assign ecchmatrix[6][418] = 1;
   assign ecchmatrix[7][418] = 1;
   assign ecchmatrix[8][418] = 0;
   assign ecchmatrix[9][418] = 1;
   assign ecchmatrix[0][419] = 1;
   assign ecchmatrix[1][419] = 1;
   assign ecchmatrix[2][419] = 0;
   assign ecchmatrix[3][419] = 1;
   assign ecchmatrix[4][419] = 0;
   assign ecchmatrix[5][419] = 1;
   assign ecchmatrix[6][419] = 1;
   assign ecchmatrix[7][419] = 0;
   assign ecchmatrix[8][419] = 1;
   assign ecchmatrix[9][419] = 1;
   assign ecchmatrix[0][420] = 1;
   assign ecchmatrix[1][420] = 1;
   assign ecchmatrix[2][420] = 0;
   assign ecchmatrix[3][420] = 1;
   assign ecchmatrix[4][420] = 0;
   assign ecchmatrix[5][420] = 1;
   assign ecchmatrix[6][420] = 0;
   assign ecchmatrix[7][420] = 1;
   assign ecchmatrix[8][420] = 1;
   assign ecchmatrix[9][420] = 1;
   assign ecchmatrix[0][421] = 1;
   assign ecchmatrix[1][421] = 1;
   assign ecchmatrix[2][421] = 0;
   assign ecchmatrix[3][421] = 1;
   assign ecchmatrix[4][421] = 0;
   assign ecchmatrix[5][421] = 0;
   assign ecchmatrix[6][421] = 1;
   assign ecchmatrix[7][421] = 1;
   assign ecchmatrix[8][421] = 1;
   assign ecchmatrix[9][421] = 1;
   assign ecchmatrix[0][422] = 1;
   assign ecchmatrix[1][422] = 1;
   assign ecchmatrix[2][422] = 0;
   assign ecchmatrix[3][422] = 0;
   assign ecchmatrix[4][422] = 1;
   assign ecchmatrix[5][422] = 1;
   assign ecchmatrix[6][422] = 1;
   assign ecchmatrix[7][422] = 1;
   assign ecchmatrix[8][422] = 1;
   assign ecchmatrix[9][422] = 0;
   assign ecchmatrix[0][423] = 1;
   assign ecchmatrix[1][423] = 1;
   assign ecchmatrix[2][423] = 0;
   assign ecchmatrix[3][423] = 0;
   assign ecchmatrix[4][423] = 1;
   assign ecchmatrix[5][423] = 1;
   assign ecchmatrix[6][423] = 1;
   assign ecchmatrix[7][423] = 1;
   assign ecchmatrix[8][423] = 0;
   assign ecchmatrix[9][423] = 1;
   assign ecchmatrix[0][424] = 1;
   assign ecchmatrix[1][424] = 1;
   assign ecchmatrix[2][424] = 0;
   assign ecchmatrix[3][424] = 0;
   assign ecchmatrix[4][424] = 1;
   assign ecchmatrix[5][424] = 1;
   assign ecchmatrix[6][424] = 1;
   assign ecchmatrix[7][424] = 0;
   assign ecchmatrix[8][424] = 1;
   assign ecchmatrix[9][424] = 1;
   assign ecchmatrix[0][425] = 1;
   assign ecchmatrix[1][425] = 1;
   assign ecchmatrix[2][425] = 0;
   assign ecchmatrix[3][425] = 0;
   assign ecchmatrix[4][425] = 1;
   assign ecchmatrix[5][425] = 1;
   assign ecchmatrix[6][425] = 0;
   assign ecchmatrix[7][425] = 1;
   assign ecchmatrix[8][425] = 1;
   assign ecchmatrix[9][425] = 1;
   assign ecchmatrix[0][426] = 1;
   assign ecchmatrix[1][426] = 1;
   assign ecchmatrix[2][426] = 0;
   assign ecchmatrix[3][426] = 0;
   assign ecchmatrix[4][426] = 1;
   assign ecchmatrix[5][426] = 0;
   assign ecchmatrix[6][426] = 1;
   assign ecchmatrix[7][426] = 1;
   assign ecchmatrix[8][426] = 1;
   assign ecchmatrix[9][426] = 1;
   assign ecchmatrix[0][427] = 1;
   assign ecchmatrix[1][427] = 1;
   assign ecchmatrix[2][427] = 0;
   assign ecchmatrix[3][427] = 0;
   assign ecchmatrix[4][427] = 0;
   assign ecchmatrix[5][427] = 1;
   assign ecchmatrix[6][427] = 1;
   assign ecchmatrix[7][427] = 1;
   assign ecchmatrix[8][427] = 1;
   assign ecchmatrix[9][427] = 1;
   assign ecchmatrix[0][428] = 1;
   assign ecchmatrix[1][428] = 0;
   assign ecchmatrix[2][428] = 1;
   assign ecchmatrix[3][428] = 1;
   assign ecchmatrix[4][428] = 1;
   assign ecchmatrix[5][428] = 1;
   assign ecchmatrix[6][428] = 1;
   assign ecchmatrix[7][428] = 1;
   assign ecchmatrix[8][428] = 0;
   assign ecchmatrix[9][428] = 0;
   assign ecchmatrix[0][429] = 1;
   assign ecchmatrix[1][429] = 0;
   assign ecchmatrix[2][429] = 1;
   assign ecchmatrix[3][429] = 1;
   assign ecchmatrix[4][429] = 1;
   assign ecchmatrix[5][429] = 1;
   assign ecchmatrix[6][429] = 1;
   assign ecchmatrix[7][429] = 0;
   assign ecchmatrix[8][429] = 1;
   assign ecchmatrix[9][429] = 0;
   assign ecchmatrix[0][430] = 1;
   assign ecchmatrix[1][430] = 0;
   assign ecchmatrix[2][430] = 1;
   assign ecchmatrix[3][430] = 1;
   assign ecchmatrix[4][430] = 1;
   assign ecchmatrix[5][430] = 1;
   assign ecchmatrix[6][430] = 1;
   assign ecchmatrix[7][430] = 0;
   assign ecchmatrix[8][430] = 0;
   assign ecchmatrix[9][430] = 1;
   assign ecchmatrix[0][431] = 1;
   assign ecchmatrix[1][431] = 0;
   assign ecchmatrix[2][431] = 1;
   assign ecchmatrix[3][431] = 1;
   assign ecchmatrix[4][431] = 1;
   assign ecchmatrix[5][431] = 1;
   assign ecchmatrix[6][431] = 0;
   assign ecchmatrix[7][431] = 1;
   assign ecchmatrix[8][431] = 1;
   assign ecchmatrix[9][431] = 0;
   assign ecchmatrix[0][432] = 1;
   assign ecchmatrix[1][432] = 0;
   assign ecchmatrix[2][432] = 1;
   assign ecchmatrix[3][432] = 1;
   assign ecchmatrix[4][432] = 1;
   assign ecchmatrix[5][432] = 1;
   assign ecchmatrix[6][432] = 0;
   assign ecchmatrix[7][432] = 1;
   assign ecchmatrix[8][432] = 0;
   assign ecchmatrix[9][432] = 1;
   assign ecchmatrix[0][433] = 1;
   assign ecchmatrix[1][433] = 0;
   assign ecchmatrix[2][433] = 1;
   assign ecchmatrix[3][433] = 1;
   assign ecchmatrix[4][433] = 1;
   assign ecchmatrix[5][433] = 1;
   assign ecchmatrix[6][433] = 0;
   assign ecchmatrix[7][433] = 0;
   assign ecchmatrix[8][433] = 1;
   assign ecchmatrix[9][433] = 1;
   assign ecchmatrix[0][434] = 1;
   assign ecchmatrix[1][434] = 0;
   assign ecchmatrix[2][434] = 1;
   assign ecchmatrix[3][434] = 1;
   assign ecchmatrix[4][434] = 1;
   assign ecchmatrix[5][434] = 0;
   assign ecchmatrix[6][434] = 1;
   assign ecchmatrix[7][434] = 1;
   assign ecchmatrix[8][434] = 1;
   assign ecchmatrix[9][434] = 0;
   assign ecchmatrix[0][435] = 1;
   assign ecchmatrix[1][435] = 0;
   assign ecchmatrix[2][435] = 1;
   assign ecchmatrix[3][435] = 1;
   assign ecchmatrix[4][435] = 1;
   assign ecchmatrix[5][435] = 0;
   assign ecchmatrix[6][435] = 1;
   assign ecchmatrix[7][435] = 1;
   assign ecchmatrix[8][435] = 0;
   assign ecchmatrix[9][435] = 1;
   assign ecchmatrix[0][436] = 1;
   assign ecchmatrix[1][436] = 0;
   assign ecchmatrix[2][436] = 1;
   assign ecchmatrix[3][436] = 1;
   assign ecchmatrix[4][436] = 1;
   assign ecchmatrix[5][436] = 0;
   assign ecchmatrix[6][436] = 1;
   assign ecchmatrix[7][436] = 0;
   assign ecchmatrix[8][436] = 1;
   assign ecchmatrix[9][436] = 1;
   assign ecchmatrix[0][437] = 1;
   assign ecchmatrix[1][437] = 0;
   assign ecchmatrix[2][437] = 1;
   assign ecchmatrix[3][437] = 1;
   assign ecchmatrix[4][437] = 1;
   assign ecchmatrix[5][437] = 0;
   assign ecchmatrix[6][437] = 0;
   assign ecchmatrix[7][437] = 1;
   assign ecchmatrix[8][437] = 1;
   assign ecchmatrix[9][437] = 1;
   assign ecchmatrix[0][438] = 1;
   assign ecchmatrix[1][438] = 0;
   assign ecchmatrix[2][438] = 1;
   assign ecchmatrix[3][438] = 1;
   assign ecchmatrix[4][438] = 0;
   assign ecchmatrix[5][438] = 1;
   assign ecchmatrix[6][438] = 1;
   assign ecchmatrix[7][438] = 1;
   assign ecchmatrix[8][438] = 1;
   assign ecchmatrix[9][438] = 0;
   assign ecchmatrix[0][439] = 1;
   assign ecchmatrix[1][439] = 0;
   assign ecchmatrix[2][439] = 1;
   assign ecchmatrix[3][439] = 1;
   assign ecchmatrix[4][439] = 0;
   assign ecchmatrix[5][439] = 1;
   assign ecchmatrix[6][439] = 1;
   assign ecchmatrix[7][439] = 1;
   assign ecchmatrix[8][439] = 0;
   assign ecchmatrix[9][439] = 1;
   assign ecchmatrix[0][440] = 1;
   assign ecchmatrix[1][440] = 0;
   assign ecchmatrix[2][440] = 1;
   assign ecchmatrix[3][440] = 1;
   assign ecchmatrix[4][440] = 0;
   assign ecchmatrix[5][440] = 1;
   assign ecchmatrix[6][440] = 1;
   assign ecchmatrix[7][440] = 0;
   assign ecchmatrix[8][440] = 1;
   assign ecchmatrix[9][440] = 1;
   assign ecchmatrix[0][441] = 1;
   assign ecchmatrix[1][441] = 0;
   assign ecchmatrix[2][441] = 1;
   assign ecchmatrix[3][441] = 1;
   assign ecchmatrix[4][441] = 0;
   assign ecchmatrix[5][441] = 1;
   assign ecchmatrix[6][441] = 0;
   assign ecchmatrix[7][441] = 1;
   assign ecchmatrix[8][441] = 1;
   assign ecchmatrix[9][441] = 1;
   assign ecchmatrix[0][442] = 1;
   assign ecchmatrix[1][442] = 0;
   assign ecchmatrix[2][442] = 1;
   assign ecchmatrix[3][442] = 1;
   assign ecchmatrix[4][442] = 0;
   assign ecchmatrix[5][442] = 0;
   assign ecchmatrix[6][442] = 1;
   assign ecchmatrix[7][442] = 1;
   assign ecchmatrix[8][442] = 1;
   assign ecchmatrix[9][442] = 1;
   assign ecchmatrix[0][443] = 1;
   assign ecchmatrix[1][443] = 0;
   assign ecchmatrix[2][443] = 1;
   assign ecchmatrix[3][443] = 0;
   assign ecchmatrix[4][443] = 1;
   assign ecchmatrix[5][443] = 1;
   assign ecchmatrix[6][443] = 1;
   assign ecchmatrix[7][443] = 1;
   assign ecchmatrix[8][443] = 1;
   assign ecchmatrix[9][443] = 0;
   assign ecchmatrix[0][444] = 1;
   assign ecchmatrix[1][444] = 0;
   assign ecchmatrix[2][444] = 1;
   assign ecchmatrix[3][444] = 0;
   assign ecchmatrix[4][444] = 1;
   assign ecchmatrix[5][444] = 1;
   assign ecchmatrix[6][444] = 1;
   assign ecchmatrix[7][444] = 1;
   assign ecchmatrix[8][444] = 0;
   assign ecchmatrix[9][444] = 1;
   assign ecchmatrix[0][445] = 1;
   assign ecchmatrix[1][445] = 0;
   assign ecchmatrix[2][445] = 1;
   assign ecchmatrix[3][445] = 0;
   assign ecchmatrix[4][445] = 1;
   assign ecchmatrix[5][445] = 1;
   assign ecchmatrix[6][445] = 1;
   assign ecchmatrix[7][445] = 0;
   assign ecchmatrix[8][445] = 1;
   assign ecchmatrix[9][445] = 1;
   assign ecchmatrix[0][446] = 1;
   assign ecchmatrix[1][446] = 0;
   assign ecchmatrix[2][446] = 1;
   assign ecchmatrix[3][446] = 0;
   assign ecchmatrix[4][446] = 1;
   assign ecchmatrix[5][446] = 1;
   assign ecchmatrix[6][446] = 0;
   assign ecchmatrix[7][446] = 1;
   assign ecchmatrix[8][446] = 1;
   assign ecchmatrix[9][446] = 1;
   assign ecchmatrix[0][447] = 1;
   assign ecchmatrix[1][447] = 0;
   assign ecchmatrix[2][447] = 1;
   assign ecchmatrix[3][447] = 0;
   assign ecchmatrix[4][447] = 1;
   assign ecchmatrix[5][447] = 0;
   assign ecchmatrix[6][447] = 1;
   assign ecchmatrix[7][447] = 1;
   assign ecchmatrix[8][447] = 1;
   assign ecchmatrix[9][447] = 1;
   assign ecchmatrix[0][448] = 1;
   assign ecchmatrix[1][448] = 0;
   assign ecchmatrix[2][448] = 1;
   assign ecchmatrix[3][448] = 0;
   assign ecchmatrix[4][448] = 0;
   assign ecchmatrix[5][448] = 1;
   assign ecchmatrix[6][448] = 1;
   assign ecchmatrix[7][448] = 1;
   assign ecchmatrix[8][448] = 1;
   assign ecchmatrix[9][448] = 1;
   assign ecchmatrix[0][449] = 1;
   assign ecchmatrix[1][449] = 0;
   assign ecchmatrix[2][449] = 0;
   assign ecchmatrix[3][449] = 1;
   assign ecchmatrix[4][449] = 1;
   assign ecchmatrix[5][449] = 1;
   assign ecchmatrix[6][449] = 1;
   assign ecchmatrix[7][449] = 1;
   assign ecchmatrix[8][449] = 1;
   assign ecchmatrix[9][449] = 0;
   assign ecchmatrix[0][450] = 1;
   assign ecchmatrix[1][450] = 0;
   assign ecchmatrix[2][450] = 0;
   assign ecchmatrix[3][450] = 1;
   assign ecchmatrix[4][450] = 1;
   assign ecchmatrix[5][450] = 1;
   assign ecchmatrix[6][450] = 1;
   assign ecchmatrix[7][450] = 1;
   assign ecchmatrix[8][450] = 0;
   assign ecchmatrix[9][450] = 1;
   assign ecchmatrix[0][451] = 1;
   assign ecchmatrix[1][451] = 0;
   assign ecchmatrix[2][451] = 0;
   assign ecchmatrix[3][451] = 1;
   assign ecchmatrix[4][451] = 1;
   assign ecchmatrix[5][451] = 1;
   assign ecchmatrix[6][451] = 1;
   assign ecchmatrix[7][451] = 0;
   assign ecchmatrix[8][451] = 1;
   assign ecchmatrix[9][451] = 1;
   assign ecchmatrix[0][452] = 1;
   assign ecchmatrix[1][452] = 0;
   assign ecchmatrix[2][452] = 0;
   assign ecchmatrix[3][452] = 1;
   assign ecchmatrix[4][452] = 1;
   assign ecchmatrix[5][452] = 1;
   assign ecchmatrix[6][452] = 0;
   assign ecchmatrix[7][452] = 1;
   assign ecchmatrix[8][452] = 1;
   assign ecchmatrix[9][452] = 1;
   assign ecchmatrix[0][453] = 1;
   assign ecchmatrix[1][453] = 0;
   assign ecchmatrix[2][453] = 0;
   assign ecchmatrix[3][453] = 1;
   assign ecchmatrix[4][453] = 1;
   assign ecchmatrix[5][453] = 0;
   assign ecchmatrix[6][453] = 1;
   assign ecchmatrix[7][453] = 1;
   assign ecchmatrix[8][453] = 1;
   assign ecchmatrix[9][453] = 1;
   assign ecchmatrix[0][454] = 1;
   assign ecchmatrix[1][454] = 0;
   assign ecchmatrix[2][454] = 0;
   assign ecchmatrix[3][454] = 1;
   assign ecchmatrix[4][454] = 0;
   assign ecchmatrix[5][454] = 1;
   assign ecchmatrix[6][454] = 1;
   assign ecchmatrix[7][454] = 1;
   assign ecchmatrix[8][454] = 1;
   assign ecchmatrix[9][454] = 1;
   assign ecchmatrix[0][455] = 1;
   assign ecchmatrix[1][455] = 0;
   assign ecchmatrix[2][455] = 0;
   assign ecchmatrix[3][455] = 0;
   assign ecchmatrix[4][455] = 1;
   assign ecchmatrix[5][455] = 1;
   assign ecchmatrix[6][455] = 1;
   assign ecchmatrix[7][455] = 1;
   assign ecchmatrix[8][455] = 1;
   assign ecchmatrix[9][455] = 1;
   assign ecchmatrix[0][456] = 0;
   assign ecchmatrix[1][456] = 1;
   assign ecchmatrix[2][456] = 1;
   assign ecchmatrix[3][456] = 1;
   assign ecchmatrix[4][456] = 1;
   assign ecchmatrix[5][456] = 1;
   assign ecchmatrix[6][456] = 1;
   assign ecchmatrix[7][456] = 1;
   assign ecchmatrix[8][456] = 0;
   assign ecchmatrix[9][456] = 0;
   assign ecchmatrix[0][457] = 0;
   assign ecchmatrix[1][457] = 1;
   assign ecchmatrix[2][457] = 1;
   assign ecchmatrix[3][457] = 1;
   assign ecchmatrix[4][457] = 1;
   assign ecchmatrix[5][457] = 1;
   assign ecchmatrix[6][457] = 1;
   assign ecchmatrix[7][457] = 0;
   assign ecchmatrix[8][457] = 1;
   assign ecchmatrix[9][457] = 0;
   assign ecchmatrix[0][458] = 0;
   assign ecchmatrix[1][458] = 1;
   assign ecchmatrix[2][458] = 1;
   assign ecchmatrix[3][458] = 1;
   assign ecchmatrix[4][458] = 1;
   assign ecchmatrix[5][458] = 1;
   assign ecchmatrix[6][458] = 1;
   assign ecchmatrix[7][458] = 0;
   assign ecchmatrix[8][458] = 0;
   assign ecchmatrix[9][458] = 1;
   assign ecchmatrix[0][459] = 0;
   assign ecchmatrix[1][459] = 1;
   assign ecchmatrix[2][459] = 1;
   assign ecchmatrix[3][459] = 1;
   assign ecchmatrix[4][459] = 1;
   assign ecchmatrix[5][459] = 1;
   assign ecchmatrix[6][459] = 0;
   assign ecchmatrix[7][459] = 1;
   assign ecchmatrix[8][459] = 1;
   assign ecchmatrix[9][459] = 0;
   assign ecchmatrix[0][460] = 0;
   assign ecchmatrix[1][460] = 1;
   assign ecchmatrix[2][460] = 1;
   assign ecchmatrix[3][460] = 1;
   assign ecchmatrix[4][460] = 1;
   assign ecchmatrix[5][460] = 1;
   assign ecchmatrix[6][460] = 0;
   assign ecchmatrix[7][460] = 1;
   assign ecchmatrix[8][460] = 0;
   assign ecchmatrix[9][460] = 1;
   assign ecchmatrix[0][461] = 0;
   assign ecchmatrix[1][461] = 1;
   assign ecchmatrix[2][461] = 1;
   assign ecchmatrix[3][461] = 1;
   assign ecchmatrix[4][461] = 1;
   assign ecchmatrix[5][461] = 1;
   assign ecchmatrix[6][461] = 0;
   assign ecchmatrix[7][461] = 0;
   assign ecchmatrix[8][461] = 1;
   assign ecchmatrix[9][461] = 1;
   assign ecchmatrix[0][462] = 0;
   assign ecchmatrix[1][462] = 1;
   assign ecchmatrix[2][462] = 1;
   assign ecchmatrix[3][462] = 1;
   assign ecchmatrix[4][462] = 1;
   assign ecchmatrix[5][462] = 0;
   assign ecchmatrix[6][462] = 1;
   assign ecchmatrix[7][462] = 1;
   assign ecchmatrix[8][462] = 1;
   assign ecchmatrix[9][462] = 0;
   assign ecchmatrix[0][463] = 0;
   assign ecchmatrix[1][463] = 1;
   assign ecchmatrix[2][463] = 1;
   assign ecchmatrix[3][463] = 1;
   assign ecchmatrix[4][463] = 1;
   assign ecchmatrix[5][463] = 0;
   assign ecchmatrix[6][463] = 1;
   assign ecchmatrix[7][463] = 1;
   assign ecchmatrix[8][463] = 0;
   assign ecchmatrix[9][463] = 1;
   assign ecchmatrix[0][464] = 0;
   assign ecchmatrix[1][464] = 1;
   assign ecchmatrix[2][464] = 1;
   assign ecchmatrix[3][464] = 1;
   assign ecchmatrix[4][464] = 1;
   assign ecchmatrix[5][464] = 0;
   assign ecchmatrix[6][464] = 1;
   assign ecchmatrix[7][464] = 0;
   assign ecchmatrix[8][464] = 1;
   assign ecchmatrix[9][464] = 1;
   assign ecchmatrix[0][465] = 0;
   assign ecchmatrix[1][465] = 1;
   assign ecchmatrix[2][465] = 1;
   assign ecchmatrix[3][465] = 1;
   assign ecchmatrix[4][465] = 1;
   assign ecchmatrix[5][465] = 0;
   assign ecchmatrix[6][465] = 0;
   assign ecchmatrix[7][465] = 1;
   assign ecchmatrix[8][465] = 1;
   assign ecchmatrix[9][465] = 1;
   assign ecchmatrix[0][466] = 0;
   assign ecchmatrix[1][466] = 1;
   assign ecchmatrix[2][466] = 1;
   assign ecchmatrix[3][466] = 1;
   assign ecchmatrix[4][466] = 0;
   assign ecchmatrix[5][466] = 1;
   assign ecchmatrix[6][466] = 1;
   assign ecchmatrix[7][466] = 1;
   assign ecchmatrix[8][466] = 1;
   assign ecchmatrix[9][466] = 0;
   assign ecchmatrix[0][467] = 0;
   assign ecchmatrix[1][467] = 1;
   assign ecchmatrix[2][467] = 1;
   assign ecchmatrix[3][467] = 1;
   assign ecchmatrix[4][467] = 0;
   assign ecchmatrix[5][467] = 1;
   assign ecchmatrix[6][467] = 1;
   assign ecchmatrix[7][467] = 1;
   assign ecchmatrix[8][467] = 0;
   assign ecchmatrix[9][467] = 1;
   assign ecchmatrix[0][468] = 0;
   assign ecchmatrix[1][468] = 1;
   assign ecchmatrix[2][468] = 1;
   assign ecchmatrix[3][468] = 1;
   assign ecchmatrix[4][468] = 0;
   assign ecchmatrix[5][468] = 1;
   assign ecchmatrix[6][468] = 1;
   assign ecchmatrix[7][468] = 0;
   assign ecchmatrix[8][468] = 1;
   assign ecchmatrix[9][468] = 1;
   assign ecchmatrix[0][469] = 0;
   assign ecchmatrix[1][469] = 1;
   assign ecchmatrix[2][469] = 1;
   assign ecchmatrix[3][469] = 1;
   assign ecchmatrix[4][469] = 0;
   assign ecchmatrix[5][469] = 1;
   assign ecchmatrix[6][469] = 0;
   assign ecchmatrix[7][469] = 1;
   assign ecchmatrix[8][469] = 1;
   assign ecchmatrix[9][469] = 1;
   assign ecchmatrix[0][470] = 0;
   assign ecchmatrix[1][470] = 1;
   assign ecchmatrix[2][470] = 1;
   assign ecchmatrix[3][470] = 1;
   assign ecchmatrix[4][470] = 0;
   assign ecchmatrix[5][470] = 0;
   assign ecchmatrix[6][470] = 1;
   assign ecchmatrix[7][470] = 1;
   assign ecchmatrix[8][470] = 1;
   assign ecchmatrix[9][470] = 1;
   assign ecchmatrix[0][471] = 0;
   assign ecchmatrix[1][471] = 1;
   assign ecchmatrix[2][471] = 1;
   assign ecchmatrix[3][471] = 0;
   assign ecchmatrix[4][471] = 1;
   assign ecchmatrix[5][471] = 1;
   assign ecchmatrix[6][471] = 1;
   assign ecchmatrix[7][471] = 1;
   assign ecchmatrix[8][471] = 1;
   assign ecchmatrix[9][471] = 0;
   assign ecchmatrix[0][472] = 0;
   assign ecchmatrix[1][472] = 1;
   assign ecchmatrix[2][472] = 1;
   assign ecchmatrix[3][472] = 0;
   assign ecchmatrix[4][472] = 1;
   assign ecchmatrix[5][472] = 1;
   assign ecchmatrix[6][472] = 1;
   assign ecchmatrix[7][472] = 1;
   assign ecchmatrix[8][472] = 0;
   assign ecchmatrix[9][472] = 1;
   assign ecchmatrix[0][473] = 0;
   assign ecchmatrix[1][473] = 1;
   assign ecchmatrix[2][473] = 1;
   assign ecchmatrix[3][473] = 0;
   assign ecchmatrix[4][473] = 1;
   assign ecchmatrix[5][473] = 1;
   assign ecchmatrix[6][473] = 1;
   assign ecchmatrix[7][473] = 0;
   assign ecchmatrix[8][473] = 1;
   assign ecchmatrix[9][473] = 1;
   assign ecchmatrix[0][474] = 0;
   assign ecchmatrix[1][474] = 1;
   assign ecchmatrix[2][474] = 1;
   assign ecchmatrix[3][474] = 0;
   assign ecchmatrix[4][474] = 1;
   assign ecchmatrix[5][474] = 1;
   assign ecchmatrix[6][474] = 0;
   assign ecchmatrix[7][474] = 1;
   assign ecchmatrix[8][474] = 1;
   assign ecchmatrix[9][474] = 1;
   assign ecchmatrix[0][475] = 0;
   assign ecchmatrix[1][475] = 1;
   assign ecchmatrix[2][475] = 1;
   assign ecchmatrix[3][475] = 0;
   assign ecchmatrix[4][475] = 1;
   assign ecchmatrix[5][475] = 0;
   assign ecchmatrix[6][475] = 1;
   assign ecchmatrix[7][475] = 1;
   assign ecchmatrix[8][475] = 1;
   assign ecchmatrix[9][475] = 1;
   assign ecchmatrix[0][476] = 0;
   assign ecchmatrix[1][476] = 1;
   assign ecchmatrix[2][476] = 1;
   assign ecchmatrix[3][476] = 0;
   assign ecchmatrix[4][476] = 0;
   assign ecchmatrix[5][476] = 1;
   assign ecchmatrix[6][476] = 1;
   assign ecchmatrix[7][476] = 1;
   assign ecchmatrix[8][476] = 1;
   assign ecchmatrix[9][476] = 1;
   assign ecchmatrix[0][477] = 0;
   assign ecchmatrix[1][477] = 1;
   assign ecchmatrix[2][477] = 0;
   assign ecchmatrix[3][477] = 1;
   assign ecchmatrix[4][477] = 1;
   assign ecchmatrix[5][477] = 1;
   assign ecchmatrix[6][477] = 1;
   assign ecchmatrix[7][477] = 1;
   assign ecchmatrix[8][477] = 1;
   assign ecchmatrix[9][477] = 0;
   assign ecchmatrix[0][478] = 0;
   assign ecchmatrix[1][478] = 1;
   assign ecchmatrix[2][478] = 0;
   assign ecchmatrix[3][478] = 1;
   assign ecchmatrix[4][478] = 1;
   assign ecchmatrix[5][478] = 1;
   assign ecchmatrix[6][478] = 1;
   assign ecchmatrix[7][478] = 1;
   assign ecchmatrix[8][478] = 0;
   assign ecchmatrix[9][478] = 1;
   assign ecchmatrix[0][479] = 0;
   assign ecchmatrix[1][479] = 1;
   assign ecchmatrix[2][479] = 0;
   assign ecchmatrix[3][479] = 1;
   assign ecchmatrix[4][479] = 1;
   assign ecchmatrix[5][479] = 1;
   assign ecchmatrix[6][479] = 1;
   assign ecchmatrix[7][479] = 0;
   assign ecchmatrix[8][479] = 1;
   assign ecchmatrix[9][479] = 1;
   assign ecchmatrix[0][480] = 0;
   assign ecchmatrix[1][480] = 1;
   assign ecchmatrix[2][480] = 0;
   assign ecchmatrix[3][480] = 1;
   assign ecchmatrix[4][480] = 1;
   assign ecchmatrix[5][480] = 1;
   assign ecchmatrix[6][480] = 0;
   assign ecchmatrix[7][480] = 1;
   assign ecchmatrix[8][480] = 1;
   assign ecchmatrix[9][480] = 1;
   assign ecchmatrix[0][481] = 0;
   assign ecchmatrix[1][481] = 1;
   assign ecchmatrix[2][481] = 0;
   assign ecchmatrix[3][481] = 1;
   assign ecchmatrix[4][481] = 1;
   assign ecchmatrix[5][481] = 0;
   assign ecchmatrix[6][481] = 1;
   assign ecchmatrix[7][481] = 1;
   assign ecchmatrix[8][481] = 1;
   assign ecchmatrix[9][481] = 1;
   assign ecchmatrix[0][482] = 0;
   assign ecchmatrix[1][482] = 1;
   assign ecchmatrix[2][482] = 0;
   assign ecchmatrix[3][482] = 1;
   assign ecchmatrix[4][482] = 0;
   assign ecchmatrix[5][482] = 1;
   assign ecchmatrix[6][482] = 1;
   assign ecchmatrix[7][482] = 1;
   assign ecchmatrix[8][482] = 1;
   assign ecchmatrix[9][482] = 1;
   assign ecchmatrix[0][483] = 0;
   assign ecchmatrix[1][483] = 1;
   assign ecchmatrix[2][483] = 0;
   assign ecchmatrix[3][483] = 0;
   assign ecchmatrix[4][483] = 1;
   assign ecchmatrix[5][483] = 1;
   assign ecchmatrix[6][483] = 1;
   assign ecchmatrix[7][483] = 1;
   assign ecchmatrix[8][483] = 1;
   assign ecchmatrix[9][483] = 1;
   assign ecchmatrix[0][484] = 0;
   assign ecchmatrix[1][484] = 0;
   assign ecchmatrix[2][484] = 1;
   assign ecchmatrix[3][484] = 1;
   assign ecchmatrix[4][484] = 1;
   assign ecchmatrix[5][484] = 1;
   assign ecchmatrix[6][484] = 1;
   assign ecchmatrix[7][484] = 1;
   assign ecchmatrix[8][484] = 1;
   assign ecchmatrix[9][484] = 0;
   assign ecchmatrix[0][485] = 0;
   assign ecchmatrix[1][485] = 0;
   assign ecchmatrix[2][485] = 1;
   assign ecchmatrix[3][485] = 1;
   assign ecchmatrix[4][485] = 1;
   assign ecchmatrix[5][485] = 1;
   assign ecchmatrix[6][485] = 1;
   assign ecchmatrix[7][485] = 1;
   assign ecchmatrix[8][485] = 0;
   assign ecchmatrix[9][485] = 1;
   assign ecchmatrix[0][486] = 0;
   assign ecchmatrix[1][486] = 0;
   assign ecchmatrix[2][486] = 1;
   assign ecchmatrix[3][486] = 1;
   assign ecchmatrix[4][486] = 1;
   assign ecchmatrix[5][486] = 1;
   assign ecchmatrix[6][486] = 1;
   assign ecchmatrix[7][486] = 0;
   assign ecchmatrix[8][486] = 1;
   assign ecchmatrix[9][486] = 1;
   assign ecchmatrix[0][487] = 0;
   assign ecchmatrix[1][487] = 0;
   assign ecchmatrix[2][487] = 1;
   assign ecchmatrix[3][487] = 1;
   assign ecchmatrix[4][487] = 1;
   assign ecchmatrix[5][487] = 1;
   assign ecchmatrix[6][487] = 0;
   assign ecchmatrix[7][487] = 1;
   assign ecchmatrix[8][487] = 1;
   assign ecchmatrix[9][487] = 1;
   assign ecchmatrix[0][488] = 0;
   assign ecchmatrix[1][488] = 0;
   assign ecchmatrix[2][488] = 1;
   assign ecchmatrix[3][488] = 1;
   assign ecchmatrix[4][488] = 1;
   assign ecchmatrix[5][488] = 0;
   assign ecchmatrix[6][488] = 1;
   assign ecchmatrix[7][488] = 1;
   assign ecchmatrix[8][488] = 1;
   assign ecchmatrix[9][488] = 1;
   assign ecchmatrix[0][489] = 0;
   assign ecchmatrix[1][489] = 0;
   assign ecchmatrix[2][489] = 1;
   assign ecchmatrix[3][489] = 1;
   assign ecchmatrix[4][489] = 0;
   assign ecchmatrix[5][489] = 1;
   assign ecchmatrix[6][489] = 1;
   assign ecchmatrix[7][489] = 1;
   assign ecchmatrix[8][489] = 1;
   assign ecchmatrix[9][489] = 1;
   assign ecchmatrix[0][490] = 0;
   assign ecchmatrix[1][490] = 0;
   assign ecchmatrix[2][490] = 1;
   assign ecchmatrix[3][490] = 0;
   assign ecchmatrix[4][490] = 1;
   assign ecchmatrix[5][490] = 1;
   assign ecchmatrix[6][490] = 1;
   assign ecchmatrix[7][490] = 1;
   assign ecchmatrix[8][490] = 1;
   assign ecchmatrix[9][490] = 1;
   assign ecchmatrix[0][491] = 0;
   assign ecchmatrix[1][491] = 0;
   assign ecchmatrix[2][491] = 0;
   assign ecchmatrix[3][491] = 1;
   assign ecchmatrix[4][491] = 1;
   assign ecchmatrix[5][491] = 1;
   assign ecchmatrix[6][491] = 1;
   assign ecchmatrix[7][491] = 1;
   assign ecchmatrix[8][491] = 1;
   assign ecchmatrix[9][491] = 1;
   assign ecchmatrix[0][492] = 1;
   assign ecchmatrix[1][492] = 1;
   assign ecchmatrix[2][492] = 1;
   assign ecchmatrix[3][492] = 1;
   assign ecchmatrix[4][492] = 1;
   assign ecchmatrix[5][492] = 1;
   assign ecchmatrix[6][492] = 1;
   assign ecchmatrix[7][492] = 1;
   assign ecchmatrix[8][492] = 1;
   assign ecchmatrix[9][492] = 0;
   assign ecchmatrix[0][493] = 1;
   assign ecchmatrix[1][493] = 1;
   assign ecchmatrix[2][493] = 1;
   assign ecchmatrix[3][493] = 1;
   assign ecchmatrix[4][493] = 1;
   assign ecchmatrix[5][493] = 1;
   assign ecchmatrix[6][493] = 1;
   assign ecchmatrix[7][493] = 1;
   assign ecchmatrix[8][493] = 0;
   assign ecchmatrix[9][493] = 1;
   assign ecchmatrix[0][494] = 1;
   assign ecchmatrix[1][494] = 1;
   assign ecchmatrix[2][494] = 1;
   assign ecchmatrix[3][494] = 1;
   assign ecchmatrix[4][494] = 1;
   assign ecchmatrix[5][494] = 1;
   assign ecchmatrix[6][494] = 1;
   assign ecchmatrix[7][494] = 0;
   assign ecchmatrix[8][494] = 1;
   assign ecchmatrix[9][494] = 1;
   assign ecchmatrix[0][495] = 1;
   assign ecchmatrix[1][495] = 1;
   assign ecchmatrix[2][495] = 1;
   assign ecchmatrix[3][495] = 1;
   assign ecchmatrix[4][495] = 1;
   assign ecchmatrix[5][495] = 1;
   assign ecchmatrix[6][495] = 0;
   assign ecchmatrix[7][495] = 1;
   assign ecchmatrix[8][495] = 1;
   assign ecchmatrix[9][495] = 1;
   assign ecchmatrix[0][496] = 1;
   assign ecchmatrix[1][496] = 1;
   assign ecchmatrix[2][496] = 1;
   assign ecchmatrix[3][496] = 1;
   assign ecchmatrix[4][496] = 1;
   assign ecchmatrix[5][496] = 0;
   assign ecchmatrix[6][496] = 1;
   assign ecchmatrix[7][496] = 1;
   assign ecchmatrix[8][496] = 1;
   assign ecchmatrix[9][496] = 1;
   assign ecchmatrix[0][497] = 1;
   assign ecchmatrix[1][497] = 1;
   assign ecchmatrix[2][497] = 1;
   assign ecchmatrix[3][497] = 1;
   assign ecchmatrix[4][497] = 0;
   assign ecchmatrix[5][497] = 1;
   assign ecchmatrix[6][497] = 1;
   assign ecchmatrix[7][497] = 1;
   assign ecchmatrix[8][497] = 1;
   assign ecchmatrix[9][497] = 1;
   assign ecchmatrix[0][498] = 1;
   assign ecchmatrix[1][498] = 1;
   assign ecchmatrix[2][498] = 1;
   assign ecchmatrix[3][498] = 0;
   assign ecchmatrix[4][498] = 1;
   assign ecchmatrix[5][498] = 1;
   assign ecchmatrix[6][498] = 1;
   assign ecchmatrix[7][498] = 1;
   assign ecchmatrix[8][498] = 1;
   assign ecchmatrix[9][498] = 1;
   assign ecchmatrix[0][499] = 1;
   assign ecchmatrix[1][499] = 1;
   assign ecchmatrix[2][499] = 0;
   assign ecchmatrix[3][499] = 1;
   assign ecchmatrix[4][499] = 1;
   assign ecchmatrix[5][499] = 1;
   assign ecchmatrix[6][499] = 1;
   assign ecchmatrix[7][499] = 1;
   assign ecchmatrix[8][499] = 1;
   assign ecchmatrix[9][499] = 1;
   assign ecchmatrix[0][500] = 1;
   assign ecchmatrix[1][500] = 0;
   assign ecchmatrix[2][500] = 1;
   assign ecchmatrix[3][500] = 1;
   assign ecchmatrix[4][500] = 1;
   assign ecchmatrix[5][500] = 1;
   assign ecchmatrix[6][500] = 1;
   assign ecchmatrix[7][500] = 1;
   assign ecchmatrix[8][500] = 1;
   assign ecchmatrix[9][500] = 1;
   assign ecchmatrix[0][501] = 0;
   assign ecchmatrix[1][501] = 1;
   assign ecchmatrix[2][501] = 1;
   assign ecchmatrix[3][501] = 1;
   assign ecchmatrix[4][501] = 1;
   assign ecchmatrix[5][501] = 1;
   assign ecchmatrix[6][501] = 1;
   assign ecchmatrix[7][501] = 1;
   assign ecchmatrix[8][501] = 1;
   assign ecchmatrix[9][501] = 1;
endmodule
