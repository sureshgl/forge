module algo_nru_1r1w (read, write, addr, din, rd_vld, rd_dout, rd_fwrd, rd_serr, rd_derr, rd_padr,
                      t1_writeA, t1_addrA, t1_dinA, t1_readB, t1_addrB, t1_doutB, t1_fwrdB, t1_serrB, t1_derrB, t1_padrB,
                      ready, clk, rst,
		              select_addr);
  
  parameter BITWDTH = 5;
  parameter WIDTH = 32;
  parameter NUMRUPT = 2;
  parameter NUMADDR = 8192;
  parameter BITADDR = 13;
  parameter NUMVROW = 1024;
  parameter BITVROW = 10;
  parameter NUMWRDS = 8;
  parameter BITWRDS = 3;
  parameter NUMPBNK = 4;     // NUMRUPT*NUMRUPT
  parameter BITPBNK = 2;
  parameter BITPADR = BITPBNK+BITADDR;
  parameter SRAM_DELAY = 2;
  parameter UPD_DELAY = 2;
  parameter FLOPIN = 0;
  parameter FLOPOUT = 0;

  input [NUMRUPT-1:0]              read;
  input [NUMRUPT-1:0]              write;
  input [NUMRUPT*BITADDR-1:0]      addr;
  input [NUMRUPT*WIDTH-1:0]        din;
  output [NUMRUPT-1:0]             rd_vld;
  output [NUMRUPT*WIDTH-1:0]       rd_dout;
  output [NUMRUPT-1:0]             rd_fwrd;
  output [NUMRUPT-1:0]             rd_serr;
  output [NUMRUPT-1:0]             rd_derr;
  output [NUMRUPT*BITPADR-1:0]     rd_padr;

  output                           ready;
  input                            clk;
  input                            rst;

  output [NUMPBNK-1:0]               t1_writeA;
  output [NUMPBNK*BITVROW-1:0]       t1_addrA;
  output [NUMPBNK*NUMWRDS*WIDTH-1:0] t1_dinA;

  output [NUMPBNK-1:0]               t1_readB;
  output [NUMPBNK*BITVROW-1:0]       t1_addrB;
  input [NUMPBNK*NUMWRDS*WIDTH-1:0]  t1_doutB;
  input [NUMPBNK-1:0]                t1_fwrdB;
  input [NUMPBNK-1:0]                t1_serrB;
  input [NUMPBNK-1:0]                t1_derrB;
  input [NUMPBNK*(BITPADR-BITPBNK-BITWRDS)-1:0] t1_padrB;

  input [BITADDR-1:0]                   select_addr;

  core_nru_1r1w #(.BITWDTH (BITWDTH), .WIDTH (WIDTH), .NUMRUPT (NUMRUPT), .NUMADDR (NUMADDR), .BITADDR (BITADDR),
                  .NUMVROW (NUMVROW), .BITVROW (BITVROW), .NUMWRDS (NUMWRDS), .BITWRDS (BITWRDS),
                  .NUMPBNK(NUMPBNK), .BITPBNK (BITPBNK), .BITPADR(BITPADR), 
                  .SRAM_DELAY (SRAM_DELAY), .UPD_DELAY (UPD_DELAY), .FLOPIN (FLOPIN), .FLOPOUT (FLOPOUT))
  core (
        .vread (read), .vwrite (write), .vaddr (addr), .vdin (din),
        .vread_vld (rd_vld), .vdout (rd_dout), .vread_fwrd (rd_fwrd), .vread_serr (rd_serr), .vread_derr (rd_derr), .vread_padr (rd_padr),
        .t1_writeA(t1_writeA), .t1_addrA(t1_addrA), .t1_dinA(t1_dinA),
        .t1_readB(t1_readB), .t1_addrB(t1_addrB), .t1_doutB(t1_doutB), .t1_fwrdB(t1_fwrdB), .t1_serrB(t1_serrB), .t1_derrB(t1_derrB), .t1_padrB(t1_padrB),
        .ready (ready), .clk (clk), .rst (rst)
        );

`ifdef FORMAL
  assume_select_addr_range: assume property (@(posedge clk) disable iff (rst) (select_addr < NUMADDR));
  assume_select_addr_stable: assume property (@(posedge clk) disable iff (rst) $stable(select_addr));

  ip_top_sva_nru_1r1w #(
                        .WIDTH       (WIDTH),
                        .BITWDTH     (BITWDTH),
                        .NUMRUPT     (NUMRUPT),
                        .NUMADDR     (NUMADDR),
                        .BITADDR     (BITADDR),
                        .NUMVROW     (NUMVROW),
                        .BITVROW     (BITVROW),
                        .NUMWRDS     (NUMWRDS),
                        .BITWRDS     (BITWRDS),
                        .NUMPBNK     (NUMPBNK),
                        .BITPBNK     (BITPBNK),
                        .BITPADR     (BITPADR),
                        .SRAM_DELAY  (SRAM_DELAY),
                        .UPD_DELAY   (UPD_DELAY),
                        .FLOPIN      (FLOPIN),
                        .FLOPOUT     (FLOPOUT))
  ip_top_sva (.*);

  ip_top_sva_2_nru_1r1w #(
                          .WIDTH       (WIDTH),
                          .NUMRUPT     (NUMRUPT),
                          .NUMADDR     (NUMADDR),
                          .BITADDR     (BITADDR),
                          .NUMVROW     (NUMVROW),
                          .BITVROW     (BITVROW),
                          .SRAM_DELAY  (SRAM_DELAY),
                          .UPD_DELAY   (UPD_DELAY))
  ip_top_sva_2 (.*);

  //`else
`elsif SIM_SVA

  genvar                                sva_int;
  generate for (sva_int=0; sva_int<WIDTH; sva_int=sva_int+1) begin : ip_top_sva
    wire [BITADDR-1:0] help_addr = sva_int;
    wire [BITWDTH-1:0] help_bit = sva_int;

    ip_top_sva_nru_1r1w #(
                          .WIDTH       (WIDTH),
                          .BITWDTH     (BITWDTH),
                          .NUMRUPT     (NUMRUPT),
                          .NUMADDR     (NUMADDR),
                          .BITADDR     (BITADDR),
                          .NUMVROW     (NUMVROW),
                          .BITVROW     (BITVROW),
                          .NUMWRDS     (NUMWRDS),
                          .BITWRDS     (BITWRDS),
                          .NUMPBNK     (NUMPBNK),
                          .BITPBNK     (BITPBNK),
                          .BITPADR     (BITPADR),
                          .SRAM_DELAY  (SRAM_DELAY),
                          .UPD_DELAY   (UPD_DELAY),
                          .FLOPIN      (FLOPIN),
                          .FLOPOUT     (FLOPOUT))
    ip_top_sva (.select_addr(help_addr), .*);
  end
  endgenerate

  ip_top_sva_2_nru_1r1w #(
                          .WIDTH       (WIDTH),
                          .NUMRUPT     (NUMRUPT),
                          .NUMADDR     (NUMADDR),
                          .BITADDR     (BITADDR),
                          .NUMVROW     (NUMVROW),
                          .BITVROW     (BITVROW),
                          .SRAM_DELAY  (SRAM_DELAY),
                          .UPD_DELAY   (UPD_DELAY))
  ip_top_sva_2 (.*);

`endif

  endmodule
