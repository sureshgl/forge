
module algo_1rfw_1rw_rl2 (clk, rst, ready,
                          write, wr_adr, din,
	                  read, rd_adr, rd_vld, rd_dout, rd_fwrd, rd_serr, rd_derr, rd_padr,
	                  t1_readA, t1_writeA, t1_addrA, t1_dinA, t1_doutA, t1_fwrdA, t1_serrA, t1_derrA, t1_padrA,
	                  t2_readA, t2_writeA, t2_addrA, t2_dinA, t2_doutA, t2_fwrdA, t2_serrA, t2_derrA, t2_padrA,
	                  t3_readA, t3_writeA, t3_addrA, t3_dinA, t3_doutA, t3_fwrdA, t3_serrA, t3_derrA, t3_padrA,
                          select_addr, select_bit);

  parameter WIDTH = 32;
  parameter BITWDTH = 5;
  parameter NUMADDR = 8192;
  parameter BITADDR = 13;
  parameter NUMVROW = 1024;
  parameter BITVROW = 10;
  parameter NUMVBNK = 8;
  parameter BITVBNK = 3;
  parameter BITPBNK = 4;
  parameter BITPADR = 14;
  parameter NUMCBNK = 2;
  parameter BITCBNK = 1;
  parameter SRAM_DELAY = 2;
  parameter FLOPIN = 0;
  parameter FLOPOUT = 0;

  input                                write;
  input [BITADDR-1:0]                  wr_adr;
  input [WIDTH-1:0]                    din;

  input                                read;
  input [BITADDR-1:0]                  rd_adr;
  output                               rd_vld;
  output [WIDTH-1:0]                   rd_dout;
  output                               rd_fwrd;
  output                               rd_serr;
  output                               rd_derr;
  output [BITPADR-1:0]                 rd_padr;

  input                                clk;
  input                                rst;
  output                               ready;

  input [BITADDR-1:0]                  select_addr;
  input [BITWDTH-1:0]                  select_bit;

  output [NUMVBNK-1:0] t1_readA;
  output [NUMVBNK-1:0] t1_writeA;
  output [NUMVBNK*BITVROW-1:0] t1_addrA;
  output [NUMVBNK*WIDTH-1:0] t1_dinA;
  input [NUMVBNK*WIDTH-1:0] t1_doutA;
  input [NUMVBNK-1:0] t1_fwrdA;
  input [NUMVBNK-1:0] t1_serrA;
  input [NUMVBNK-1:0] t1_derrA;
  input [NUMVBNK*(BITPADR-BITPBNK)-1:0] t1_padrA;

  output [NUMCBNK-1:0] t2_readA;
  output [NUMCBNK-1:0] t2_writeA;
  output [NUMCBNK*BITVROW-1:0] t2_addrA;
  output [NUMCBNK*WIDTH-1:0] t2_dinA;
  input [NUMCBNK*WIDTH-1:0] t2_doutA;
  input [NUMCBNK-1:0] t2_fwrdA;
  input [NUMCBNK-1:0] t2_serrA;
  input [NUMCBNK-1:0] t2_derrA;
  input [NUMCBNK*(BITPADR-BITPBNK)-1:0] t2_padrA;

  output [NUMCBNK-1:0] t3_readA;
  output [NUMCBNK-1:0] t3_writeA;
  output [NUMCBNK*BITVROW-1:0] t3_addrA;
  output [NUMCBNK*(BITVBNK+1)-1:0] t3_dinA;
  input [NUMCBNK*(BITVBNK+1)-1:0] t3_doutA;
  input [NUMCBNK-1:0] t3_fwrdA;
  input [NUMCBNK-1:0] t3_serrA;
  input [NUMCBNK-1:0] t3_derrA;
  input [NUMCBNK*(BITPADR-BITPBNK)-1:0] t3_padrA;

  core_1rfw_1rw_rl2 #(.WIDTH (WIDTH), .BITWDTH (BITWDTH), .NUMADDR (NUMADDR), .BITADDR (BITADDR),
                      .NUMVROW (NUMVROW), .BITVROW (BITVROW), .NUMVBNK (NUMVBNK), .BITVBNK (BITVBNK), .BITPBNK (BITPBNK), .BITPADR (BITPADR),
                      .NUMCBNK (NUMCBNK), .BITCBNK (BITCBNK),
                      .SRAM_DELAY (SRAM_DELAY), .FLOPIN (FLOPIN), .FLOPOUT (FLOPOUT))
    core (.vread (read), .vrdaddr (rd_adr), .vread_vld (rd_vld), .vdout (rd_dout),
          .vread_fwrd (rd_fwrd), .vread_serr (rd_serr), .vread_derr (rd_derr), .vread_padr (rd_padr),
          .vwrite (write), .vwraddr (wr_adr), .vdin (din),
          .t1_readA(t1_readA), .t1_writeA(t1_writeA), .t1_addrA(t1_addrA), .t1_dinA(t1_dinA), .t1_doutA(t1_doutA),
          .t1_fwrdA(t1_fwrdA), .t1_serrA(t1_serrA), .t1_derrA(t1_derrA), .t1_padrA(t1_padrA),
          .t2_readA(t2_readA), .t2_writeA(t2_writeA), .t2_addrA(t2_addrA), .t2_dinA(t2_dinA), .t2_doutA(t2_doutA),
          .t2_fwrdA(t2_fwrdA), .t2_serrA(t2_serrA), .t2_derrA(t2_derrA), .t2_padrA(t2_padrA),
          .t3_readA(t3_readA), .t3_writeA(t3_writeA), .t3_addrA(t3_addrA), .t3_dinA(t3_dinA), .t3_doutA(t3_doutA),
          .t3_fwrdA(t3_fwrdA), .t3_serrA(t3_serrA), .t3_derrA(t3_derrA), .t3_padrA(t3_padrA),
          .ready (ready), .clk (clk), .rst (rst),
          .select_addr (select_addr), .select_bit (select_bit));

`ifdef FORMAL
assume_select_addr_range: assume property (@(posedge clk) disable iff (rst) (select_addr < NUMADDR));
assume_select_addr_stable: assume property (@(posedge clk) disable iff (rst) $stable(select_addr));
assume_select_bit_range: assume property (@(posedge clk) disable iff (rst) (select_bit < WIDTH));
assume_select_bit_stable: assume property (@(posedge clk) disable iff (rst) $stable(select_bit));

ip_top_sva_1rfw_1rw_rl2 #(
     .WIDTH       (WIDTH),
     .BITWDTH     (BITWDTH),
     .NUMADDR     (NUMADDR),
     .BITADDR     (BITADDR),
     .NUMVROW     (NUMVROW),
     .BITVROW     (BITVROW),
     .NUMVBNK     (NUMVBNK),
     .BITVBNK     (BITVBNK),
     .BITPBNK     (BITPBNK),
     .BITPADR     (BITPADR),
     .NUMCBNK     (NUMCBNK),
     .BITCBNK     (BITCBNK),
     .SRAM_DELAY  (SRAM_DELAY),
     .FLOPIN      (FLOPIN),
     .FLOPOUT     (FLOPOUT))
ip_top_sva (.*);

ip_top_sva_2_1rfw_1rw_rl2 #(
     .WIDTH       (WIDTH),
     .BITWDTH     (BITWDTH),
     .NUMADDR     (NUMADDR),
     .BITADDR     (BITADDR),
     .NUMVROW     (NUMVROW),
     .BITVROW     (BITVROW),
     .NUMVBNK     (NUMVBNK),
     .BITVBNK     (BITVBNK),
     .NUMCBNK     (NUMCBNK),
     .BITCBNK     (BITCBNK),
     .SRAM_DELAY  (SRAM_DELAY))
ip_top_sva_2 (.*);

`elsif SIM_SVA

genvar sva_int;
generate for (sva_int=0; sva_int<1; sva_int=sva_int+1) begin
  wire [BITADDR-1:0] help_addr = sva_int;
  wire [BITWDTH-1:0] help_bit = sva_int;
ip_top_sva_1rfw_1rw_rl2 #(
     .WIDTH       (WIDTH),
     .BITWDTH     (BITWDTH),
     .NUMADDR     (NUMADDR),
     .BITADDR     (BITADDR),
     .NUMVROW     (NUMVROW),
     .BITVROW     (BITVROW),
     .NUMVBNK     (NUMVBNK),
     .BITVBNK     (BITVBNK),
     .BITPBNK     (BITPBNK),
     .BITPADR     (BITPADR),
     .NUMCBNK     (NUMCBNK),
     .BITCBNK     (BITCBNK),
     .SRAM_DELAY  (SRAM_DELAY),
     .FLOPIN      (FLOPIN),
     .FLOPOUT     (FLOPOUT))
ip_top_sva (.select_addr(help_addr), .select_bit (help_bit), .*);
end
endgenerate

ip_top_sva_2_1rfw_1rw_rl2 #(
     .WIDTH       (WIDTH),
     .BITWDTH     (BITWDTH),
     .NUMADDR     (NUMADDR),
     .BITADDR     (BITADDR),
     .NUMVROW     (NUMVROW),
     .BITVROW     (BITVROW),
     .NUMVBNK     (NUMVBNK),
     .BITVBNK     (BITVBNK),
     .NUMCBNK     (NUMCBNK),
     .BITCBNK     (BITCBNK),
     .SRAM_DELAY  (SRAM_DELAY))
ip_top_sva_2 (.*);

`endif

endmodule
