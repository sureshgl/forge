module ip_top_sva_afifo (

                         );

  parameter WIDTH   = 32;
  parameter NUMWRDS = 16;
  parameter BITAPTR =  8;
  parameter BITWRDS = 4;

endmodule // ip_top_sva_afifo

module ip_top_sva_2_afifo (

                         );

  parameter WIDTH   = 32;
  parameter NUMWRDS = 16;
  parameter BITAPTR =  8;
  parameter BITWRDS = 4;

endmodule // ip_top_sva_afifo
