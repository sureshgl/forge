`define ARB_FIFO_PKT_THRESHOLD_OFFSET	32'h0
`define ARB_FIFO_PKT_THRESHOLD_SIZE	16
`define ARB_FIFO_PKT_THRESHOLD_SIZE_IN_WORDS	1

`define ARB_FIFO_PKT_THRESHOLD_THRESH_SIZE	16
`define ARB_FIFO_PKT_THRESHOLD_THRESH_START_OFFSET	0
`define ARB_FIFO_PKT_THRESHOLD_THRESH_RANGE	[15:0]
`define ARB_FIFO_PKT_THRESHOLD_THRESH_RST_VALUE	16'hF0'h16'hF0




`define PROC_PKT_THRESHOLD_0_OFFSET	32'h8
`define PROC_PKT_THRESHOLD_0_SIZE	33
`define PROC_PKT_THRESHOLD_0_SIZE_IN_WORDS	6
`define PROC_PKT_THRESHOLD_1_OFFSET	32'ha
`define PROC_PKT_THRESHOLD_1_SIZE	33
`define PROC_PKT_THRESHOLD_1_SIZE_IN_WORDS	6
`define PROC_PKT_THRESHOLD_2_OFFSET	32'hc
`define PROC_PKT_THRESHOLD_2_SIZE	33
`define PROC_PKT_THRESHOLD_2_SIZE_IN_WORDS	6

`define PROC_PKT_THRESHOLD_THRESH_SIZE	33
`define PROC_PKT_THRESHOLD_THRESH_START_OFFSET	0
`define PROC_PKT_THRESHOLD_THRESH_RANGE	[32:0]
`define PROC_PKT_THRESHOLD_THRESH_RST_VALUE	16'h0FF'h16'h0FF




`define DUMMYREG_OFFSET	32'h10
`define DUMMYREG_SIZE	39
`define DUMMYREG_SIZE_IN_WORDS	2

`define DUMMYREG_THRESH_SIZE	39
`define DUMMYREG_THRESH_START_OFFSET	0
`define DUMMYREG_THRESH_RANGE	[38:0]
`define DUMMYREG_THRESH_RST_VALUE	16'hF0'h16'hF0




`define DUMMY_REG_0_OFFSET	32'h20
`define DUMMY_REG_0_SIZE	65
`define DUMMY_REG_0_SIZE_IN_WORDS	18
`define DUMMY_REG_1_OFFSET	32'h23
`define DUMMY_REG_1_SIZE	65
`define DUMMY_REG_1_SIZE_IN_WORDS	18
`define DUMMY_REG_2_OFFSET	32'h26
`define DUMMY_REG_2_SIZE	65
`define DUMMY_REG_2_SIZE_IN_WORDS	18
`define DUMMY_REG_3_OFFSET	32'h29
`define DUMMY_REG_3_SIZE	65
`define DUMMY_REG_3_SIZE_IN_WORDS	18
`define DUMMY_REG_4_OFFSET	32'h2c
`define DUMMY_REG_4_SIZE	65
`define DUMMY_REG_4_SIZE_IN_WORDS	18
`define DUMMY_REG_5_OFFSET	32'h2f
`define DUMMY_REG_5_SIZE	65
`define DUMMY_REG_5_SIZE_IN_WORDS	18

`define DUMMY_REG_THRESH_SIZE	65
`define DUMMY_REG_THRESH_START_OFFSET	0
`define DUMMY_REG_THRESH_RANGE	[64:0]
`define DUMMY_REG_THRESH_RST_VALUE	16'h0FF'h16'h0FF




`define MEM_1_OFFSET	32'h40
`define MEM_1_NUMROWS	32
`define MEM_1_WIDTH	16
`define MEM_1_WIDTH_IN_WORDS	1

`define MEM_1_FL1_SIZE	11
`define MEM_1_FL1_START_OFFSET	0
`define MEM_1_FL1_RANGE	[10:0]
`define MEM_1_FL1_RST_VALUE	0'h0




`define MEM_2_0_OFFSET	32'h80
`define MEM_2_0_NUMROWS	32
`define MEM_2_0_WIDTH	64
`define MEM_2_0_WIDTH_IN_WORDS	2
`define MEM_2_1_OFFSET	32'hc0
`define MEM_2_1_NUMROWS	32
`define MEM_2_1_WIDTH	64
`define MEM_2_1_WIDTH_IN_WORDS	2
`define MEM_2_2_OFFSET	32'h100
`define MEM_2_2_NUMROWS	32
`define MEM_2_2_WIDTH	64
`define MEM_2_2_WIDTH_IN_WORDS	2

`define MEM_2_FL1_SIZE	13
`define MEM_2_FL1_START_OFFSET	0
`define MEM_2_FL1_RANGE	[12:0]
`define MEM_2_FL1_RST_VALUE	0'h0




`define MEM_3_OFFSET	32'h200
`define MEM_3_NUMROWS	128
`define MEM_3_WIDTH	64
`define MEM_3_WIDTH_IN_WORDS	2

`define MEM_3_FL1_SIZE	14
`define MEM_3_FL1_START_OFFSET	0
`define MEM_3_FL1_RANGE	[13:0]
`define MEM_3_FL1_RST_VALUE	0'h0





