//////////////////////////////////////////////////////////////////////////////
// Copyright 2010, Cisco Systems, Inc.
// All Rights Reserved. 
// 
// This is UNPUBLISHED PROPRIETARY SOURCE CODE of Cisco Systems, Inc; 
// the contents of this file may not be disclosed to third parties, copied or 
// duplicated in any form, in whole or in part, without the prior written 
// permission of Cisco Systems, Inc. 
// 
// RESTRICTED RIGHTS LEGEND: 
// Use, duplication or disclosure by the Government is subject to restrictions 
// as set forth in subdivision (c)(1)(ii) of the Rights in Technical Data 
// and Computer Software clause at DFARS 252.227-7013, and/or in similar or 
// successor clauses in the FAR, DOD or NASA FAR Supplement. Unpublished - 
// rights reserved under the Copyright Laws of the United States. 
//
//////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
//This file is auto-generated using rdlWrapGen.pl
//
//Do not modify this file modify the Source file (RDL).
//Filename = IpfBlock0RdlWrapCepDefines.vh.

 `ifndef  __IPF_BLOCK0_RDL_WRAP_CEP_DEFINES_VH_
 `define  __IPF_BLOCK0_RDL_WRAP_CEP_DEFINES_VH_
 `include "MemRdlCommStructs.vh"


 `define IPF_LINK_LIST_MMR0_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR0_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR0_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR0_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR0_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR1_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR1_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR1_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR1_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR1_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR10_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR10_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR10_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR10_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR10_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR11_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR11_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR11_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR11_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR11_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR12_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR12_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR12_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR12_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR12_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR13_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR13_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR13_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR13_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR13_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR14_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR14_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR14_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR14_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR14_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR15_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR15_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR15_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR15_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR15_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR16_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR16_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR16_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR16_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR16_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR17_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR17_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR17_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR17_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR17_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR18_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR18_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR18_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR18_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR18_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR19_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR19_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR19_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR19_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR19_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR2_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR2_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR2_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR2_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR2_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR3_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR3_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR3_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR3_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR3_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR4_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR4_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR4_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR4_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR4_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR5_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR5_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR5_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR5_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR5_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR6_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR6_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR6_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR6_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR6_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR7_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR7_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR7_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR7_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR7_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR8_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR8_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR8_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR8_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR8_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)

 `define IPF_LINK_LIST_MMR9_RDLTOMEM_TYPE RdlToMemCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR9_MEMTORDL_TYPE MemToRdlCpuEccFulleBus_t

 `define IPF_LINK_LIST_MMR9_CEP_PARAM .RDL_TO_MEM_BUS_TYPE	(`IPF_LINK_LIST_MMR9_RDLTOMEM_TYPE), \
 .MEM_TO_RDL_BUS_TYPE	(`IPF_LINK_LIST_MMR9_MEMTORDL_TYPE) \
, .CPU	(1), .ECC	(1), .PARITY	(0), .BIP	(0), .ELAM	(1), .ELAM_HAS_DOUT	(1)


//Depth 
`define IPFLINKLISTMMR0_NUM                                            512
`define IPFLINKLISTMMR1_NUM                                            512
`define IPFLINKLISTMMR2_NUM                                            512
`define IPFLINKLISTMMR3_NUM                                            512
`define IPFLINKLISTMMR4_NUM                                            512
`define IPFLINKLISTMMR5_NUM                                            512
`define IPFLINKLISTMMR6_NUM                                            512
`define IPFLINKLISTMMR7_NUM                                            512
`define IPFLINKLISTMMR8_NUM                                            512
`define IPFLINKLISTMMR9_NUM                                            512
`define IPFLINKLISTMMR10_NUM                                           512
`define IPFLINKLISTMMR11_NUM                                           512
`define IPFLINKLISTMMR12_NUM                                           512
`define IPFLINKLISTMMR13_NUM                                           512
`define IPFLINKLISTMMR14_NUM                                           512
`define IPFLINKLISTMMR15_NUM                                           512
`define IPFLINKLISTMMR16_NUM                                           512
`define IPFLINKLISTMMR17_NUM                                           512
`define IPFLINKLISTMMR18_NUM                                           1024
`define IPFLINKLISTMMR19_NUM                                           1024
//Physical width
`define IPFLINKLISTMMR0_PHY_WIDTH                                        16
`define IPFLINKLISTMMR1_PHY_WIDTH                                        16
`define IPFLINKLISTMMR2_PHY_WIDTH                                        16
`define IPFLINKLISTMMR3_PHY_WIDTH                                        16
`define IPFLINKLISTMMR4_PHY_WIDTH                                        16
`define IPFLINKLISTMMR5_PHY_WIDTH                                        16
`define IPFLINKLISTMMR6_PHY_WIDTH                                        10
`define IPFLINKLISTMMR7_PHY_WIDTH                                        10
`define IPFLINKLISTMMR8_PHY_WIDTH                                        10
`define IPFLINKLISTMMR9_PHY_WIDTH                                       568
`define IPFLINKLISTMMR10_PHY_WIDTH                                      568
`define IPFLINKLISTMMR11_PHY_WIDTH                                      568
`define IPFLINKLISTMMR12_PHY_WIDTH                                      568
`define IPFLINKLISTMMR13_PHY_WIDTH                                      568
`define IPFLINKLISTMMR14_PHY_WIDTH                                      568
`define IPFLINKLISTMMR15_PHY_WIDTH                                       10
`define IPFLINKLISTMMR16_PHY_WIDTH                                       10
`define IPFLINKLISTMMR17_PHY_WIDTH                                       10
`define IPFLINKLISTMMR18_PHY_WIDTH                                       11
`define IPFLINKLISTMMR19_PHY_WIDTH                                       11
//Logical width
`define IPFLINKLISTMMR0_WIDTH                                            32
`define IPFLINKLISTMMR1_WIDTH                                            32
`define IPFLINKLISTMMR2_WIDTH                                            32
`define IPFLINKLISTMMR3_WIDTH                                            32
`define IPFLINKLISTMMR4_WIDTH                                            32
`define IPFLINKLISTMMR5_WIDTH                                            32
`define IPFLINKLISTMMR6_WIDTH                                            32
`define IPFLINKLISTMMR7_WIDTH                                            32
`define IPFLINKLISTMMR8_WIDTH                                            32
`define IPFLINKLISTMMR9_WIDTH                                          1024
`define IPFLINKLISTMMR10_WIDTH                                         1024
`define IPFLINKLISTMMR11_WIDTH                                         1024
`define IPFLINKLISTMMR12_WIDTH                                         1024
`define IPFLINKLISTMMR13_WIDTH                                         1024
`define IPFLINKLISTMMR14_WIDTH                                         1024
`define IPFLINKLISTMMR15_WIDTH                                           32
`define IPFLINKLISTMMR16_WIDTH                                           32
`define IPFLINKLISTMMR17_WIDTH                                           32
`define IPFLINKLISTMMR18_WIDTH                                           32
`define IPFLINKLISTMMR19_WIDTH                                           32
//Logical mask
`define IPFLINKLISTMMR0_MASK           32'b11111111111111110000000000000000
`define IPFLINKLISTMMR1_MASK           32'b11111111111111110000000000000000
`define IPFLINKLISTMMR2_MASK           32'b11111111111111110000000000000000
`define IPFLINKLISTMMR3_MASK           32'b11111111111111110000000000000000
`define IPFLINKLISTMMR4_MASK           32'b11111111111111110000000000000000
`define IPFLINKLISTMMR5_MASK           32'b11111111111111110000000000000000
`define IPFLINKLISTMMR6_MASK           32'b11111111111111111111110000000000
`define IPFLINKLISTMMR7_MASK           32'b11111111111111111111110000000000
`define IPFLINKLISTMMR8_MASK           32'b11111111111111111111110000000000
`define IPFLINKLISTMMR9_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define IPFLINKLISTMMR10_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define IPFLINKLISTMMR11_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define IPFLINKLISTMMR12_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define IPFLINKLISTMMR13_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define IPFLINKLISTMMR14_MASK 1024'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
`define IPFLINKLISTMMR15_MASK          32'b11111111111111111111110000000000
`define IPFLINKLISTMMR16_MASK          32'b11111111111111111111110000000000
`define IPFLINKLISTMMR17_MASK          32'b11111111111111111111110000000000
`define IPFLINKLISTMMR18_MASK          32'b11111111111111111111100000000000
`define IPFLINKLISTMMR19_MASK          32'b11111111111111111111100000000000

 `endif
